`define FPGA_BUILD 1
`include "alu_definitions.v"
`include "decode_definitions.v"
`include "issue_definitions.v"
`include "lsu_definitions.v"
`include "global_definitions.v"
module decoder_10_to_1024 (out,in);
  output [1023:0] out;
  input [9:0] in;
// %%start_veriperl
// my $i;
// for($i=0; $i<1024; $i=$i+1)
// {
//   print "  assign out[$i] = (in == 10'd$i) ? 1'b1 : 1'b0;\n";
// }
// %%stop_veriperl
  assign out[0] = (in == 10'd0) ? 1'b1 : 1'b0;
  assign out[1] = (in == 10'd1) ? 1'b1 : 1'b0;
  assign out[2] = (in == 10'd2) ? 1'b1 : 1'b0;
  assign out[3] = (in == 10'd3) ? 1'b1 : 1'b0;
  assign out[4] = (in == 10'd4) ? 1'b1 : 1'b0;
  assign out[5] = (in == 10'd5) ? 1'b1 : 1'b0;
  assign out[6] = (in == 10'd6) ? 1'b1 : 1'b0;
  assign out[7] = (in == 10'd7) ? 1'b1 : 1'b0;
  assign out[8] = (in == 10'd8) ? 1'b1 : 1'b0;
  assign out[9] = (in == 10'd9) ? 1'b1 : 1'b0;
  assign out[10] = (in == 10'd10) ? 1'b1 : 1'b0;
  assign out[11] = (in == 10'd11) ? 1'b1 : 1'b0;
  assign out[12] = (in == 10'd12) ? 1'b1 : 1'b0;
  assign out[13] = (in == 10'd13) ? 1'b1 : 1'b0;
  assign out[14] = (in == 10'd14) ? 1'b1 : 1'b0;
  assign out[15] = (in == 10'd15) ? 1'b1 : 1'b0;
  assign out[16] = (in == 10'd16) ? 1'b1 : 1'b0;
  assign out[17] = (in == 10'd17) ? 1'b1 : 1'b0;
  assign out[18] = (in == 10'd18) ? 1'b1 : 1'b0;
  assign out[19] = (in == 10'd19) ? 1'b1 : 1'b0;
  assign out[20] = (in == 10'd20) ? 1'b1 : 1'b0;
  assign out[21] = (in == 10'd21) ? 1'b1 : 1'b0;
  assign out[22] = (in == 10'd22) ? 1'b1 : 1'b0;
  assign out[23] = (in == 10'd23) ? 1'b1 : 1'b0;
  assign out[24] = (in == 10'd24) ? 1'b1 : 1'b0;
  assign out[25] = (in == 10'd25) ? 1'b1 : 1'b0;
  assign out[26] = (in == 10'd26) ? 1'b1 : 1'b0;
  assign out[27] = (in == 10'd27) ? 1'b1 : 1'b0;
  assign out[28] = (in == 10'd28) ? 1'b1 : 1'b0;
  assign out[29] = (in == 10'd29) ? 1'b1 : 1'b0;
  assign out[30] = (in == 10'd30) ? 1'b1 : 1'b0;
  assign out[31] = (in == 10'd31) ? 1'b1 : 1'b0;
  assign out[32] = (in == 10'd32) ? 1'b1 : 1'b0;
  assign out[33] = (in == 10'd33) ? 1'b1 : 1'b0;
  assign out[34] = (in == 10'd34) ? 1'b1 : 1'b0;
  assign out[35] = (in == 10'd35) ? 1'b1 : 1'b0;
  assign out[36] = (in == 10'd36) ? 1'b1 : 1'b0;
  assign out[37] = (in == 10'd37) ? 1'b1 : 1'b0;
  assign out[38] = (in == 10'd38) ? 1'b1 : 1'b0;
  assign out[39] = (in == 10'd39) ? 1'b1 : 1'b0;
  assign out[40] = (in == 10'd40) ? 1'b1 : 1'b0;
  assign out[41] = (in == 10'd41) ? 1'b1 : 1'b0;
  assign out[42] = (in == 10'd42) ? 1'b1 : 1'b0;
  assign out[43] = (in == 10'd43) ? 1'b1 : 1'b0;
  assign out[44] = (in == 10'd44) ? 1'b1 : 1'b0;
  assign out[45] = (in == 10'd45) ? 1'b1 : 1'b0;
  assign out[46] = (in == 10'd46) ? 1'b1 : 1'b0;
  assign out[47] = (in == 10'd47) ? 1'b1 : 1'b0;
  assign out[48] = (in == 10'd48) ? 1'b1 : 1'b0;
  assign out[49] = (in == 10'd49) ? 1'b1 : 1'b0;
  assign out[50] = (in == 10'd50) ? 1'b1 : 1'b0;
  assign out[51] = (in == 10'd51) ? 1'b1 : 1'b0;
  assign out[52] = (in == 10'd52) ? 1'b1 : 1'b0;
  assign out[53] = (in == 10'd53) ? 1'b1 : 1'b0;
  assign out[54] = (in == 10'd54) ? 1'b1 : 1'b0;
  assign out[55] = (in == 10'd55) ? 1'b1 : 1'b0;
  assign out[56] = (in == 10'd56) ? 1'b1 : 1'b0;
  assign out[57] = (in == 10'd57) ? 1'b1 : 1'b0;
  assign out[58] = (in == 10'd58) ? 1'b1 : 1'b0;
  assign out[59] = (in == 10'd59) ? 1'b1 : 1'b0;
  assign out[60] = (in == 10'd60) ? 1'b1 : 1'b0;
  assign out[61] = (in == 10'd61) ? 1'b1 : 1'b0;
  assign out[62] = (in == 10'd62) ? 1'b1 : 1'b0;
  assign out[63] = (in == 10'd63) ? 1'b1 : 1'b0;
  assign out[64] = (in == 10'd64) ? 1'b1 : 1'b0;
  assign out[65] = (in == 10'd65) ? 1'b1 : 1'b0;
  assign out[66] = (in == 10'd66) ? 1'b1 : 1'b0;
  assign out[67] = (in == 10'd67) ? 1'b1 : 1'b0;
  assign out[68] = (in == 10'd68) ? 1'b1 : 1'b0;
  assign out[69] = (in == 10'd69) ? 1'b1 : 1'b0;
  assign out[70] = (in == 10'd70) ? 1'b1 : 1'b0;
  assign out[71] = (in == 10'd71) ? 1'b1 : 1'b0;
  assign out[72] = (in == 10'd72) ? 1'b1 : 1'b0;
  assign out[73] = (in == 10'd73) ? 1'b1 : 1'b0;
  assign out[74] = (in == 10'd74) ? 1'b1 : 1'b0;
  assign out[75] = (in == 10'd75) ? 1'b1 : 1'b0;
  assign out[76] = (in == 10'd76) ? 1'b1 : 1'b0;
  assign out[77] = (in == 10'd77) ? 1'b1 : 1'b0;
  assign out[78] = (in == 10'd78) ? 1'b1 : 1'b0;
  assign out[79] = (in == 10'd79) ? 1'b1 : 1'b0;
  assign out[80] = (in == 10'd80) ? 1'b1 : 1'b0;
  assign out[81] = (in == 10'd81) ? 1'b1 : 1'b0;
  assign out[82] = (in == 10'd82) ? 1'b1 : 1'b0;
  assign out[83] = (in == 10'd83) ? 1'b1 : 1'b0;
  assign out[84] = (in == 10'd84) ? 1'b1 : 1'b0;
  assign out[85] = (in == 10'd85) ? 1'b1 : 1'b0;
  assign out[86] = (in == 10'd86) ? 1'b1 : 1'b0;
  assign out[87] = (in == 10'd87) ? 1'b1 : 1'b0;
  assign out[88] = (in == 10'd88) ? 1'b1 : 1'b0;
  assign out[89] = (in == 10'd89) ? 1'b1 : 1'b0;
  assign out[90] = (in == 10'd90) ? 1'b1 : 1'b0;
  assign out[91] = (in == 10'd91) ? 1'b1 : 1'b0;
  assign out[92] = (in == 10'd92) ? 1'b1 : 1'b0;
  assign out[93] = (in == 10'd93) ? 1'b1 : 1'b0;
  assign out[94] = (in == 10'd94) ? 1'b1 : 1'b0;
  assign out[95] = (in == 10'd95) ? 1'b1 : 1'b0;
  assign out[96] = (in == 10'd96) ? 1'b1 : 1'b0;
  assign out[97] = (in == 10'd97) ? 1'b1 : 1'b0;
  assign out[98] = (in == 10'd98) ? 1'b1 : 1'b0;
  assign out[99] = (in == 10'd99) ? 1'b1 : 1'b0;
  assign out[100] = (in == 10'd100) ? 1'b1 : 1'b0;
  assign out[101] = (in == 10'd101) ? 1'b1 : 1'b0;
  assign out[102] = (in == 10'd102) ? 1'b1 : 1'b0;
  assign out[103] = (in == 10'd103) ? 1'b1 : 1'b0;
  assign out[104] = (in == 10'd104) ? 1'b1 : 1'b0;
  assign out[105] = (in == 10'd105) ? 1'b1 : 1'b0;
  assign out[106] = (in == 10'd106) ? 1'b1 : 1'b0;
  assign out[107] = (in == 10'd107) ? 1'b1 : 1'b0;
  assign out[108] = (in == 10'd108) ? 1'b1 : 1'b0;
  assign out[109] = (in == 10'd109) ? 1'b1 : 1'b0;
  assign out[110] = (in == 10'd110) ? 1'b1 : 1'b0;
  assign out[111] = (in == 10'd111) ? 1'b1 : 1'b0;
  assign out[112] = (in == 10'd112) ? 1'b1 : 1'b0;
  assign out[113] = (in == 10'd113) ? 1'b1 : 1'b0;
  assign out[114] = (in == 10'd114) ? 1'b1 : 1'b0;
  assign out[115] = (in == 10'd115) ? 1'b1 : 1'b0;
  assign out[116] = (in == 10'd116) ? 1'b1 : 1'b0;
  assign out[117] = (in == 10'd117) ? 1'b1 : 1'b0;
  assign out[118] = (in == 10'd118) ? 1'b1 : 1'b0;
  assign out[119] = (in == 10'd119) ? 1'b1 : 1'b0;
  assign out[120] = (in == 10'd120) ? 1'b1 : 1'b0;
  assign out[121] = (in == 10'd121) ? 1'b1 : 1'b0;
  assign out[122] = (in == 10'd122) ? 1'b1 : 1'b0;
  assign out[123] = (in == 10'd123) ? 1'b1 : 1'b0;
  assign out[124] = (in == 10'd124) ? 1'b1 : 1'b0;
  assign out[125] = (in == 10'd125) ? 1'b1 : 1'b0;
  assign out[126] = (in == 10'd126) ? 1'b1 : 1'b0;
  assign out[127] = (in == 10'd127) ? 1'b1 : 1'b0;
  assign out[128] = (in == 10'd128) ? 1'b1 : 1'b0;
  assign out[129] = (in == 10'd129) ? 1'b1 : 1'b0;
  assign out[130] = (in == 10'd130) ? 1'b1 : 1'b0;
  assign out[131] = (in == 10'd131) ? 1'b1 : 1'b0;
  assign out[132] = (in == 10'd132) ? 1'b1 : 1'b0;
  assign out[133] = (in == 10'd133) ? 1'b1 : 1'b0;
  assign out[134] = (in == 10'd134) ? 1'b1 : 1'b0;
  assign out[135] = (in == 10'd135) ? 1'b1 : 1'b0;
  assign out[136] = (in == 10'd136) ? 1'b1 : 1'b0;
  assign out[137] = (in == 10'd137) ? 1'b1 : 1'b0;
  assign out[138] = (in == 10'd138) ? 1'b1 : 1'b0;
  assign out[139] = (in == 10'd139) ? 1'b1 : 1'b0;
  assign out[140] = (in == 10'd140) ? 1'b1 : 1'b0;
  assign out[141] = (in == 10'd141) ? 1'b1 : 1'b0;
  assign out[142] = (in == 10'd142) ? 1'b1 : 1'b0;
  assign out[143] = (in == 10'd143) ? 1'b1 : 1'b0;
  assign out[144] = (in == 10'd144) ? 1'b1 : 1'b0;
  assign out[145] = (in == 10'd145) ? 1'b1 : 1'b0;
  assign out[146] = (in == 10'd146) ? 1'b1 : 1'b0;
  assign out[147] = (in == 10'd147) ? 1'b1 : 1'b0;
  assign out[148] = (in == 10'd148) ? 1'b1 : 1'b0;
  assign out[149] = (in == 10'd149) ? 1'b1 : 1'b0;
  assign out[150] = (in == 10'd150) ? 1'b1 : 1'b0;
  assign out[151] = (in == 10'd151) ? 1'b1 : 1'b0;
  assign out[152] = (in == 10'd152) ? 1'b1 : 1'b0;
  assign out[153] = (in == 10'd153) ? 1'b1 : 1'b0;
  assign out[154] = (in == 10'd154) ? 1'b1 : 1'b0;
  assign out[155] = (in == 10'd155) ? 1'b1 : 1'b0;
  assign out[156] = (in == 10'd156) ? 1'b1 : 1'b0;
  assign out[157] = (in == 10'd157) ? 1'b1 : 1'b0;
  assign out[158] = (in == 10'd158) ? 1'b1 : 1'b0;
  assign out[159] = (in == 10'd159) ? 1'b1 : 1'b0;
  assign out[160] = (in == 10'd160) ? 1'b1 : 1'b0;
  assign out[161] = (in == 10'd161) ? 1'b1 : 1'b0;
  assign out[162] = (in == 10'd162) ? 1'b1 : 1'b0;
  assign out[163] = (in == 10'd163) ? 1'b1 : 1'b0;
  assign out[164] = (in == 10'd164) ? 1'b1 : 1'b0;
  assign out[165] = (in == 10'd165) ? 1'b1 : 1'b0;
  assign out[166] = (in == 10'd166) ? 1'b1 : 1'b0;
  assign out[167] = (in == 10'd167) ? 1'b1 : 1'b0;
  assign out[168] = (in == 10'd168) ? 1'b1 : 1'b0;
  assign out[169] = (in == 10'd169) ? 1'b1 : 1'b0;
  assign out[170] = (in == 10'd170) ? 1'b1 : 1'b0;
  assign out[171] = (in == 10'd171) ? 1'b1 : 1'b0;
  assign out[172] = (in == 10'd172) ? 1'b1 : 1'b0;
  assign out[173] = (in == 10'd173) ? 1'b1 : 1'b0;
  assign out[174] = (in == 10'd174) ? 1'b1 : 1'b0;
  assign out[175] = (in == 10'd175) ? 1'b1 : 1'b0;
  assign out[176] = (in == 10'd176) ? 1'b1 : 1'b0;
  assign out[177] = (in == 10'd177) ? 1'b1 : 1'b0;
  assign out[178] = (in == 10'd178) ? 1'b1 : 1'b0;
  assign out[179] = (in == 10'd179) ? 1'b1 : 1'b0;
  assign out[180] = (in == 10'd180) ? 1'b1 : 1'b0;
  assign out[181] = (in == 10'd181) ? 1'b1 : 1'b0;
  assign out[182] = (in == 10'd182) ? 1'b1 : 1'b0;
  assign out[183] = (in == 10'd183) ? 1'b1 : 1'b0;
  assign out[184] = (in == 10'd184) ? 1'b1 : 1'b0;
  assign out[185] = (in == 10'd185) ? 1'b1 : 1'b0;
  assign out[186] = (in == 10'd186) ? 1'b1 : 1'b0;
  assign out[187] = (in == 10'd187) ? 1'b1 : 1'b0;
  assign out[188] = (in == 10'd188) ? 1'b1 : 1'b0;
  assign out[189] = (in == 10'd189) ? 1'b1 : 1'b0;
  assign out[190] = (in == 10'd190) ? 1'b1 : 1'b0;
  assign out[191] = (in == 10'd191) ? 1'b1 : 1'b0;
  assign out[192] = (in == 10'd192) ? 1'b1 : 1'b0;
  assign out[193] = (in == 10'd193) ? 1'b1 : 1'b0;
  assign out[194] = (in == 10'd194) ? 1'b1 : 1'b0;
  assign out[195] = (in == 10'd195) ? 1'b1 : 1'b0;
  assign out[196] = (in == 10'd196) ? 1'b1 : 1'b0;
  assign out[197] = (in == 10'd197) ? 1'b1 : 1'b0;
  assign out[198] = (in == 10'd198) ? 1'b1 : 1'b0;
  assign out[199] = (in == 10'd199) ? 1'b1 : 1'b0;
  assign out[200] = (in == 10'd200) ? 1'b1 : 1'b0;
  assign out[201] = (in == 10'd201) ? 1'b1 : 1'b0;
  assign out[202] = (in == 10'd202) ? 1'b1 : 1'b0;
  assign out[203] = (in == 10'd203) ? 1'b1 : 1'b0;
  assign out[204] = (in == 10'd204) ? 1'b1 : 1'b0;
  assign out[205] = (in == 10'd205) ? 1'b1 : 1'b0;
  assign out[206] = (in == 10'd206) ? 1'b1 : 1'b0;
  assign out[207] = (in == 10'd207) ? 1'b1 : 1'b0;
  assign out[208] = (in == 10'd208) ? 1'b1 : 1'b0;
  assign out[209] = (in == 10'd209) ? 1'b1 : 1'b0;
  assign out[210] = (in == 10'd210) ? 1'b1 : 1'b0;
  assign out[211] = (in == 10'd211) ? 1'b1 : 1'b0;
  assign out[212] = (in == 10'd212) ? 1'b1 : 1'b0;
  assign out[213] = (in == 10'd213) ? 1'b1 : 1'b0;
  assign out[214] = (in == 10'd214) ? 1'b1 : 1'b0;
  assign out[215] = (in == 10'd215) ? 1'b1 : 1'b0;
  assign out[216] = (in == 10'd216) ? 1'b1 : 1'b0;
  assign out[217] = (in == 10'd217) ? 1'b1 : 1'b0;
  assign out[218] = (in == 10'd218) ? 1'b1 : 1'b0;
  assign out[219] = (in == 10'd219) ? 1'b1 : 1'b0;
  assign out[220] = (in == 10'd220) ? 1'b1 : 1'b0;
  assign out[221] = (in == 10'd221) ? 1'b1 : 1'b0;
  assign out[222] = (in == 10'd222) ? 1'b1 : 1'b0;
  assign out[223] = (in == 10'd223) ? 1'b1 : 1'b0;
  assign out[224] = (in == 10'd224) ? 1'b1 : 1'b0;
  assign out[225] = (in == 10'd225) ? 1'b1 : 1'b0;
  assign out[226] = (in == 10'd226) ? 1'b1 : 1'b0;
  assign out[227] = (in == 10'd227) ? 1'b1 : 1'b0;
  assign out[228] = (in == 10'd228) ? 1'b1 : 1'b0;
  assign out[229] = (in == 10'd229) ? 1'b1 : 1'b0;
  assign out[230] = (in == 10'd230) ? 1'b1 : 1'b0;
  assign out[231] = (in == 10'd231) ? 1'b1 : 1'b0;
  assign out[232] = (in == 10'd232) ? 1'b1 : 1'b0;
  assign out[233] = (in == 10'd233) ? 1'b1 : 1'b0;
  assign out[234] = (in == 10'd234) ? 1'b1 : 1'b0;
  assign out[235] = (in == 10'd235) ? 1'b1 : 1'b0;
  assign out[236] = (in == 10'd236) ? 1'b1 : 1'b0;
  assign out[237] = (in == 10'd237) ? 1'b1 : 1'b0;
  assign out[238] = (in == 10'd238) ? 1'b1 : 1'b0;
  assign out[239] = (in == 10'd239) ? 1'b1 : 1'b0;
  assign out[240] = (in == 10'd240) ? 1'b1 : 1'b0;
  assign out[241] = (in == 10'd241) ? 1'b1 : 1'b0;
  assign out[242] = (in == 10'd242) ? 1'b1 : 1'b0;
  assign out[243] = (in == 10'd243) ? 1'b1 : 1'b0;
  assign out[244] = (in == 10'd244) ? 1'b1 : 1'b0;
  assign out[245] = (in == 10'd245) ? 1'b1 : 1'b0;
  assign out[246] = (in == 10'd246) ? 1'b1 : 1'b0;
  assign out[247] = (in == 10'd247) ? 1'b1 : 1'b0;
  assign out[248] = (in == 10'd248) ? 1'b1 : 1'b0;
  assign out[249] = (in == 10'd249) ? 1'b1 : 1'b0;
  assign out[250] = (in == 10'd250) ? 1'b1 : 1'b0;
  assign out[251] = (in == 10'd251) ? 1'b1 : 1'b0;
  assign out[252] = (in == 10'd252) ? 1'b1 : 1'b0;
  assign out[253] = (in == 10'd253) ? 1'b1 : 1'b0;
  assign out[254] = (in == 10'd254) ? 1'b1 : 1'b0;
  assign out[255] = (in == 10'd255) ? 1'b1 : 1'b0;
  assign out[256] = (in == 10'd256) ? 1'b1 : 1'b0;
  assign out[257] = (in == 10'd257) ? 1'b1 : 1'b0;
  assign out[258] = (in == 10'd258) ? 1'b1 : 1'b0;
  assign out[259] = (in == 10'd259) ? 1'b1 : 1'b0;
  assign out[260] = (in == 10'd260) ? 1'b1 : 1'b0;
  assign out[261] = (in == 10'd261) ? 1'b1 : 1'b0;
  assign out[262] = (in == 10'd262) ? 1'b1 : 1'b0;
  assign out[263] = (in == 10'd263) ? 1'b1 : 1'b0;
  assign out[264] = (in == 10'd264) ? 1'b1 : 1'b0;
  assign out[265] = (in == 10'd265) ? 1'b1 : 1'b0;
  assign out[266] = (in == 10'd266) ? 1'b1 : 1'b0;
  assign out[267] = (in == 10'd267) ? 1'b1 : 1'b0;
  assign out[268] = (in == 10'd268) ? 1'b1 : 1'b0;
  assign out[269] = (in == 10'd269) ? 1'b1 : 1'b0;
  assign out[270] = (in == 10'd270) ? 1'b1 : 1'b0;
  assign out[271] = (in == 10'd271) ? 1'b1 : 1'b0;
  assign out[272] = (in == 10'd272) ? 1'b1 : 1'b0;
  assign out[273] = (in == 10'd273) ? 1'b1 : 1'b0;
  assign out[274] = (in == 10'd274) ? 1'b1 : 1'b0;
  assign out[275] = (in == 10'd275) ? 1'b1 : 1'b0;
  assign out[276] = (in == 10'd276) ? 1'b1 : 1'b0;
  assign out[277] = (in == 10'd277) ? 1'b1 : 1'b0;
  assign out[278] = (in == 10'd278) ? 1'b1 : 1'b0;
  assign out[279] = (in == 10'd279) ? 1'b1 : 1'b0;
  assign out[280] = (in == 10'd280) ? 1'b1 : 1'b0;
  assign out[281] = (in == 10'd281) ? 1'b1 : 1'b0;
  assign out[282] = (in == 10'd282) ? 1'b1 : 1'b0;
  assign out[283] = (in == 10'd283) ? 1'b1 : 1'b0;
  assign out[284] = (in == 10'd284) ? 1'b1 : 1'b0;
  assign out[285] = (in == 10'd285) ? 1'b1 : 1'b0;
  assign out[286] = (in == 10'd286) ? 1'b1 : 1'b0;
  assign out[287] = (in == 10'd287) ? 1'b1 : 1'b0;
  assign out[288] = (in == 10'd288) ? 1'b1 : 1'b0;
  assign out[289] = (in == 10'd289) ? 1'b1 : 1'b0;
  assign out[290] = (in == 10'd290) ? 1'b1 : 1'b0;
  assign out[291] = (in == 10'd291) ? 1'b1 : 1'b0;
  assign out[292] = (in == 10'd292) ? 1'b1 : 1'b0;
  assign out[293] = (in == 10'd293) ? 1'b1 : 1'b0;
  assign out[294] = (in == 10'd294) ? 1'b1 : 1'b0;
  assign out[295] = (in == 10'd295) ? 1'b1 : 1'b0;
  assign out[296] = (in == 10'd296) ? 1'b1 : 1'b0;
  assign out[297] = (in == 10'd297) ? 1'b1 : 1'b0;
  assign out[298] = (in == 10'd298) ? 1'b1 : 1'b0;
  assign out[299] = (in == 10'd299) ? 1'b1 : 1'b0;
  assign out[300] = (in == 10'd300) ? 1'b1 : 1'b0;
  assign out[301] = (in == 10'd301) ? 1'b1 : 1'b0;
  assign out[302] = (in == 10'd302) ? 1'b1 : 1'b0;
  assign out[303] = (in == 10'd303) ? 1'b1 : 1'b0;
  assign out[304] = (in == 10'd304) ? 1'b1 : 1'b0;
  assign out[305] = (in == 10'd305) ? 1'b1 : 1'b0;
  assign out[306] = (in == 10'd306) ? 1'b1 : 1'b0;
  assign out[307] = (in == 10'd307) ? 1'b1 : 1'b0;
  assign out[308] = (in == 10'd308) ? 1'b1 : 1'b0;
  assign out[309] = (in == 10'd309) ? 1'b1 : 1'b0;
  assign out[310] = (in == 10'd310) ? 1'b1 : 1'b0;
  assign out[311] = (in == 10'd311) ? 1'b1 : 1'b0;
  assign out[312] = (in == 10'd312) ? 1'b1 : 1'b0;
  assign out[313] = (in == 10'd313) ? 1'b1 : 1'b0;
  assign out[314] = (in == 10'd314) ? 1'b1 : 1'b0;
  assign out[315] = (in == 10'd315) ? 1'b1 : 1'b0;
  assign out[316] = (in == 10'd316) ? 1'b1 : 1'b0;
  assign out[317] = (in == 10'd317) ? 1'b1 : 1'b0;
  assign out[318] = (in == 10'd318) ? 1'b1 : 1'b0;
  assign out[319] = (in == 10'd319) ? 1'b1 : 1'b0;
  assign out[320] = (in == 10'd320) ? 1'b1 : 1'b0;
  assign out[321] = (in == 10'd321) ? 1'b1 : 1'b0;
  assign out[322] = (in == 10'd322) ? 1'b1 : 1'b0;
  assign out[323] = (in == 10'd323) ? 1'b1 : 1'b0;
  assign out[324] = (in == 10'd324) ? 1'b1 : 1'b0;
  assign out[325] = (in == 10'd325) ? 1'b1 : 1'b0;
  assign out[326] = (in == 10'd326) ? 1'b1 : 1'b0;
  assign out[327] = (in == 10'd327) ? 1'b1 : 1'b0;
  assign out[328] = (in == 10'd328) ? 1'b1 : 1'b0;
  assign out[329] = (in == 10'd329) ? 1'b1 : 1'b0;
  assign out[330] = (in == 10'd330) ? 1'b1 : 1'b0;
  assign out[331] = (in == 10'd331) ? 1'b1 : 1'b0;
  assign out[332] = (in == 10'd332) ? 1'b1 : 1'b0;
  assign out[333] = (in == 10'd333) ? 1'b1 : 1'b0;
  assign out[334] = (in == 10'd334) ? 1'b1 : 1'b0;
  assign out[335] = (in == 10'd335) ? 1'b1 : 1'b0;
  assign out[336] = (in == 10'd336) ? 1'b1 : 1'b0;
  assign out[337] = (in == 10'd337) ? 1'b1 : 1'b0;
  assign out[338] = (in == 10'd338) ? 1'b1 : 1'b0;
  assign out[339] = (in == 10'd339) ? 1'b1 : 1'b0;
  assign out[340] = (in == 10'd340) ? 1'b1 : 1'b0;
  assign out[341] = (in == 10'd341) ? 1'b1 : 1'b0;
  assign out[342] = (in == 10'd342) ? 1'b1 : 1'b0;
  assign out[343] = (in == 10'd343) ? 1'b1 : 1'b0;
  assign out[344] = (in == 10'd344) ? 1'b1 : 1'b0;
  assign out[345] = (in == 10'd345) ? 1'b1 : 1'b0;
  assign out[346] = (in == 10'd346) ? 1'b1 : 1'b0;
  assign out[347] = (in == 10'd347) ? 1'b1 : 1'b0;
  assign out[348] = (in == 10'd348) ? 1'b1 : 1'b0;
  assign out[349] = (in == 10'd349) ? 1'b1 : 1'b0;
  assign out[350] = (in == 10'd350) ? 1'b1 : 1'b0;
  assign out[351] = (in == 10'd351) ? 1'b1 : 1'b0;
  assign out[352] = (in == 10'd352) ? 1'b1 : 1'b0;
  assign out[353] = (in == 10'd353) ? 1'b1 : 1'b0;
  assign out[354] = (in == 10'd354) ? 1'b1 : 1'b0;
  assign out[355] = (in == 10'd355) ? 1'b1 : 1'b0;
  assign out[356] = (in == 10'd356) ? 1'b1 : 1'b0;
  assign out[357] = (in == 10'd357) ? 1'b1 : 1'b0;
  assign out[358] = (in == 10'd358) ? 1'b1 : 1'b0;
  assign out[359] = (in == 10'd359) ? 1'b1 : 1'b0;
  assign out[360] = (in == 10'd360) ? 1'b1 : 1'b0;
  assign out[361] = (in == 10'd361) ? 1'b1 : 1'b0;
  assign out[362] = (in == 10'd362) ? 1'b1 : 1'b0;
  assign out[363] = (in == 10'd363) ? 1'b1 : 1'b0;
  assign out[364] = (in == 10'd364) ? 1'b1 : 1'b0;
  assign out[365] = (in == 10'd365) ? 1'b1 : 1'b0;
  assign out[366] = (in == 10'd366) ? 1'b1 : 1'b0;
  assign out[367] = (in == 10'd367) ? 1'b1 : 1'b0;
  assign out[368] = (in == 10'd368) ? 1'b1 : 1'b0;
  assign out[369] = (in == 10'd369) ? 1'b1 : 1'b0;
  assign out[370] = (in == 10'd370) ? 1'b1 : 1'b0;
  assign out[371] = (in == 10'd371) ? 1'b1 : 1'b0;
  assign out[372] = (in == 10'd372) ? 1'b1 : 1'b0;
  assign out[373] = (in == 10'd373) ? 1'b1 : 1'b0;
  assign out[374] = (in == 10'd374) ? 1'b1 : 1'b0;
  assign out[375] = (in == 10'd375) ? 1'b1 : 1'b0;
  assign out[376] = (in == 10'd376) ? 1'b1 : 1'b0;
  assign out[377] = (in == 10'd377) ? 1'b1 : 1'b0;
  assign out[378] = (in == 10'd378) ? 1'b1 : 1'b0;
  assign out[379] = (in == 10'd379) ? 1'b1 : 1'b0;
  assign out[380] = (in == 10'd380) ? 1'b1 : 1'b0;
  assign out[381] = (in == 10'd381) ? 1'b1 : 1'b0;
  assign out[382] = (in == 10'd382) ? 1'b1 : 1'b0;
  assign out[383] = (in == 10'd383) ? 1'b1 : 1'b0;
  assign out[384] = (in == 10'd384) ? 1'b1 : 1'b0;
  assign out[385] = (in == 10'd385) ? 1'b1 : 1'b0;
  assign out[386] = (in == 10'd386) ? 1'b1 : 1'b0;
  assign out[387] = (in == 10'd387) ? 1'b1 : 1'b0;
  assign out[388] = (in == 10'd388) ? 1'b1 : 1'b0;
  assign out[389] = (in == 10'd389) ? 1'b1 : 1'b0;
  assign out[390] = (in == 10'd390) ? 1'b1 : 1'b0;
  assign out[391] = (in == 10'd391) ? 1'b1 : 1'b0;
  assign out[392] = (in == 10'd392) ? 1'b1 : 1'b0;
  assign out[393] = (in == 10'd393) ? 1'b1 : 1'b0;
  assign out[394] = (in == 10'd394) ? 1'b1 : 1'b0;
  assign out[395] = (in == 10'd395) ? 1'b1 : 1'b0;
  assign out[396] = (in == 10'd396) ? 1'b1 : 1'b0;
  assign out[397] = (in == 10'd397) ? 1'b1 : 1'b0;
  assign out[398] = (in == 10'd398) ? 1'b1 : 1'b0;
  assign out[399] = (in == 10'd399) ? 1'b1 : 1'b0;
  assign out[400] = (in == 10'd400) ? 1'b1 : 1'b0;
  assign out[401] = (in == 10'd401) ? 1'b1 : 1'b0;
  assign out[402] = (in == 10'd402) ? 1'b1 : 1'b0;
  assign out[403] = (in == 10'd403) ? 1'b1 : 1'b0;
  assign out[404] = (in == 10'd404) ? 1'b1 : 1'b0;
  assign out[405] = (in == 10'd405) ? 1'b1 : 1'b0;
  assign out[406] = (in == 10'd406) ? 1'b1 : 1'b0;
  assign out[407] = (in == 10'd407) ? 1'b1 : 1'b0;
  assign out[408] = (in == 10'd408) ? 1'b1 : 1'b0;
  assign out[409] = (in == 10'd409) ? 1'b1 : 1'b0;
  assign out[410] = (in == 10'd410) ? 1'b1 : 1'b0;
  assign out[411] = (in == 10'd411) ? 1'b1 : 1'b0;
  assign out[412] = (in == 10'd412) ? 1'b1 : 1'b0;
  assign out[413] = (in == 10'd413) ? 1'b1 : 1'b0;
  assign out[414] = (in == 10'd414) ? 1'b1 : 1'b0;
  assign out[415] = (in == 10'd415) ? 1'b1 : 1'b0;
  assign out[416] = (in == 10'd416) ? 1'b1 : 1'b0;
  assign out[417] = (in == 10'd417) ? 1'b1 : 1'b0;
  assign out[418] = (in == 10'd418) ? 1'b1 : 1'b0;
  assign out[419] = (in == 10'd419) ? 1'b1 : 1'b0;
  assign out[420] = (in == 10'd420) ? 1'b1 : 1'b0;
  assign out[421] = (in == 10'd421) ? 1'b1 : 1'b0;
  assign out[422] = (in == 10'd422) ? 1'b1 : 1'b0;
  assign out[423] = (in == 10'd423) ? 1'b1 : 1'b0;
  assign out[424] = (in == 10'd424) ? 1'b1 : 1'b0;
  assign out[425] = (in == 10'd425) ? 1'b1 : 1'b0;
  assign out[426] = (in == 10'd426) ? 1'b1 : 1'b0;
  assign out[427] = (in == 10'd427) ? 1'b1 : 1'b0;
  assign out[428] = (in == 10'd428) ? 1'b1 : 1'b0;
  assign out[429] = (in == 10'd429) ? 1'b1 : 1'b0;
  assign out[430] = (in == 10'd430) ? 1'b1 : 1'b0;
  assign out[431] = (in == 10'd431) ? 1'b1 : 1'b0;
  assign out[432] = (in == 10'd432) ? 1'b1 : 1'b0;
  assign out[433] = (in == 10'd433) ? 1'b1 : 1'b0;
  assign out[434] = (in == 10'd434) ? 1'b1 : 1'b0;
  assign out[435] = (in == 10'd435) ? 1'b1 : 1'b0;
  assign out[436] = (in == 10'd436) ? 1'b1 : 1'b0;
  assign out[437] = (in == 10'd437) ? 1'b1 : 1'b0;
  assign out[438] = (in == 10'd438) ? 1'b1 : 1'b0;
  assign out[439] = (in == 10'd439) ? 1'b1 : 1'b0;
  assign out[440] = (in == 10'd440) ? 1'b1 : 1'b0;
  assign out[441] = (in == 10'd441) ? 1'b1 : 1'b0;
  assign out[442] = (in == 10'd442) ? 1'b1 : 1'b0;
  assign out[443] = (in == 10'd443) ? 1'b1 : 1'b0;
  assign out[444] = (in == 10'd444) ? 1'b1 : 1'b0;
  assign out[445] = (in == 10'd445) ? 1'b1 : 1'b0;
  assign out[446] = (in == 10'd446) ? 1'b1 : 1'b0;
  assign out[447] = (in == 10'd447) ? 1'b1 : 1'b0;
  assign out[448] = (in == 10'd448) ? 1'b1 : 1'b0;
  assign out[449] = (in == 10'd449) ? 1'b1 : 1'b0;
  assign out[450] = (in == 10'd450) ? 1'b1 : 1'b0;
  assign out[451] = (in == 10'd451) ? 1'b1 : 1'b0;
  assign out[452] = (in == 10'd452) ? 1'b1 : 1'b0;
  assign out[453] = (in == 10'd453) ? 1'b1 : 1'b0;
  assign out[454] = (in == 10'd454) ? 1'b1 : 1'b0;
  assign out[455] = (in == 10'd455) ? 1'b1 : 1'b0;
  assign out[456] = (in == 10'd456) ? 1'b1 : 1'b0;
  assign out[457] = (in == 10'd457) ? 1'b1 : 1'b0;
  assign out[458] = (in == 10'd458) ? 1'b1 : 1'b0;
  assign out[459] = (in == 10'd459) ? 1'b1 : 1'b0;
  assign out[460] = (in == 10'd460) ? 1'b1 : 1'b0;
  assign out[461] = (in == 10'd461) ? 1'b1 : 1'b0;
  assign out[462] = (in == 10'd462) ? 1'b1 : 1'b0;
  assign out[463] = (in == 10'd463) ? 1'b1 : 1'b0;
  assign out[464] = (in == 10'd464) ? 1'b1 : 1'b0;
  assign out[465] = (in == 10'd465) ? 1'b1 : 1'b0;
  assign out[466] = (in == 10'd466) ? 1'b1 : 1'b0;
  assign out[467] = (in == 10'd467) ? 1'b1 : 1'b0;
  assign out[468] = (in == 10'd468) ? 1'b1 : 1'b0;
  assign out[469] = (in == 10'd469) ? 1'b1 : 1'b0;
  assign out[470] = (in == 10'd470) ? 1'b1 : 1'b0;
  assign out[471] = (in == 10'd471) ? 1'b1 : 1'b0;
  assign out[472] = (in == 10'd472) ? 1'b1 : 1'b0;
  assign out[473] = (in == 10'd473) ? 1'b1 : 1'b0;
  assign out[474] = (in == 10'd474) ? 1'b1 : 1'b0;
  assign out[475] = (in == 10'd475) ? 1'b1 : 1'b0;
  assign out[476] = (in == 10'd476) ? 1'b1 : 1'b0;
  assign out[477] = (in == 10'd477) ? 1'b1 : 1'b0;
  assign out[478] = (in == 10'd478) ? 1'b1 : 1'b0;
  assign out[479] = (in == 10'd479) ? 1'b1 : 1'b0;
  assign out[480] = (in == 10'd480) ? 1'b1 : 1'b0;
  assign out[481] = (in == 10'd481) ? 1'b1 : 1'b0;
  assign out[482] = (in == 10'd482) ? 1'b1 : 1'b0;
  assign out[483] = (in == 10'd483) ? 1'b1 : 1'b0;
  assign out[484] = (in == 10'd484) ? 1'b1 : 1'b0;
  assign out[485] = (in == 10'd485) ? 1'b1 : 1'b0;
  assign out[486] = (in == 10'd486) ? 1'b1 : 1'b0;
  assign out[487] = (in == 10'd487) ? 1'b1 : 1'b0;
  assign out[488] = (in == 10'd488) ? 1'b1 : 1'b0;
  assign out[489] = (in == 10'd489) ? 1'b1 : 1'b0;
  assign out[490] = (in == 10'd490) ? 1'b1 : 1'b0;
  assign out[491] = (in == 10'd491) ? 1'b1 : 1'b0;
  assign out[492] = (in == 10'd492) ? 1'b1 : 1'b0;
  assign out[493] = (in == 10'd493) ? 1'b1 : 1'b0;
  assign out[494] = (in == 10'd494) ? 1'b1 : 1'b0;
  assign out[495] = (in == 10'd495) ? 1'b1 : 1'b0;
  assign out[496] = (in == 10'd496) ? 1'b1 : 1'b0;
  assign out[497] = (in == 10'd497) ? 1'b1 : 1'b0;
  assign out[498] = (in == 10'd498) ? 1'b1 : 1'b0;
  assign out[499] = (in == 10'd499) ? 1'b1 : 1'b0;
  assign out[500] = (in == 10'd500) ? 1'b1 : 1'b0;
  assign out[501] = (in == 10'd501) ? 1'b1 : 1'b0;
  assign out[502] = (in == 10'd502) ? 1'b1 : 1'b0;
  assign out[503] = (in == 10'd503) ? 1'b1 : 1'b0;
  assign out[504] = (in == 10'd504) ? 1'b1 : 1'b0;
  assign out[505] = (in == 10'd505) ? 1'b1 : 1'b0;
  assign out[506] = (in == 10'd506) ? 1'b1 : 1'b0;
  assign out[507] = (in == 10'd507) ? 1'b1 : 1'b0;
  assign out[508] = (in == 10'd508) ? 1'b1 : 1'b0;
  assign out[509] = (in == 10'd509) ? 1'b1 : 1'b0;
  assign out[510] = (in == 10'd510) ? 1'b1 : 1'b0;
  assign out[511] = (in == 10'd511) ? 1'b1 : 1'b0;
  assign out[512] = (in == 10'd512) ? 1'b1 : 1'b0;
  assign out[513] = (in == 10'd513) ? 1'b1 : 1'b0;
  assign out[514] = (in == 10'd514) ? 1'b1 : 1'b0;
  assign out[515] = (in == 10'd515) ? 1'b1 : 1'b0;
  assign out[516] = (in == 10'd516) ? 1'b1 : 1'b0;
  assign out[517] = (in == 10'd517) ? 1'b1 : 1'b0;
  assign out[518] = (in == 10'd518) ? 1'b1 : 1'b0;
  assign out[519] = (in == 10'd519) ? 1'b1 : 1'b0;
  assign out[520] = (in == 10'd520) ? 1'b1 : 1'b0;
  assign out[521] = (in == 10'd521) ? 1'b1 : 1'b0;
  assign out[522] = (in == 10'd522) ? 1'b1 : 1'b0;
  assign out[523] = (in == 10'd523) ? 1'b1 : 1'b0;
  assign out[524] = (in == 10'd524) ? 1'b1 : 1'b0;
  assign out[525] = (in == 10'd525) ? 1'b1 : 1'b0;
  assign out[526] = (in == 10'd526) ? 1'b1 : 1'b0;
  assign out[527] = (in == 10'd527) ? 1'b1 : 1'b0;
  assign out[528] = (in == 10'd528) ? 1'b1 : 1'b0;
  assign out[529] = (in == 10'd529) ? 1'b1 : 1'b0;
  assign out[530] = (in == 10'd530) ? 1'b1 : 1'b0;
  assign out[531] = (in == 10'd531) ? 1'b1 : 1'b0;
  assign out[532] = (in == 10'd532) ? 1'b1 : 1'b0;
  assign out[533] = (in == 10'd533) ? 1'b1 : 1'b0;
  assign out[534] = (in == 10'd534) ? 1'b1 : 1'b0;
  assign out[535] = (in == 10'd535) ? 1'b1 : 1'b0;
  assign out[536] = (in == 10'd536) ? 1'b1 : 1'b0;
  assign out[537] = (in == 10'd537) ? 1'b1 : 1'b0;
  assign out[538] = (in == 10'd538) ? 1'b1 : 1'b0;
  assign out[539] = (in == 10'd539) ? 1'b1 : 1'b0;
  assign out[540] = (in == 10'd540) ? 1'b1 : 1'b0;
  assign out[541] = (in == 10'd541) ? 1'b1 : 1'b0;
  assign out[542] = (in == 10'd542) ? 1'b1 : 1'b0;
  assign out[543] = (in == 10'd543) ? 1'b1 : 1'b0;
  assign out[544] = (in == 10'd544) ? 1'b1 : 1'b0;
  assign out[545] = (in == 10'd545) ? 1'b1 : 1'b0;
  assign out[546] = (in == 10'd546) ? 1'b1 : 1'b0;
  assign out[547] = (in == 10'd547) ? 1'b1 : 1'b0;
  assign out[548] = (in == 10'd548) ? 1'b1 : 1'b0;
  assign out[549] = (in == 10'd549) ? 1'b1 : 1'b0;
  assign out[550] = (in == 10'd550) ? 1'b1 : 1'b0;
  assign out[551] = (in == 10'd551) ? 1'b1 : 1'b0;
  assign out[552] = (in == 10'd552) ? 1'b1 : 1'b0;
  assign out[553] = (in == 10'd553) ? 1'b1 : 1'b0;
  assign out[554] = (in == 10'd554) ? 1'b1 : 1'b0;
  assign out[555] = (in == 10'd555) ? 1'b1 : 1'b0;
  assign out[556] = (in == 10'd556) ? 1'b1 : 1'b0;
  assign out[557] = (in == 10'd557) ? 1'b1 : 1'b0;
  assign out[558] = (in == 10'd558) ? 1'b1 : 1'b0;
  assign out[559] = (in == 10'd559) ? 1'b1 : 1'b0;
  assign out[560] = (in == 10'd560) ? 1'b1 : 1'b0;
  assign out[561] = (in == 10'd561) ? 1'b1 : 1'b0;
  assign out[562] = (in == 10'd562) ? 1'b1 : 1'b0;
  assign out[563] = (in == 10'd563) ? 1'b1 : 1'b0;
  assign out[564] = (in == 10'd564) ? 1'b1 : 1'b0;
  assign out[565] = (in == 10'd565) ? 1'b1 : 1'b0;
  assign out[566] = (in == 10'd566) ? 1'b1 : 1'b0;
  assign out[567] = (in == 10'd567) ? 1'b1 : 1'b0;
  assign out[568] = (in == 10'd568) ? 1'b1 : 1'b0;
  assign out[569] = (in == 10'd569) ? 1'b1 : 1'b0;
  assign out[570] = (in == 10'd570) ? 1'b1 : 1'b0;
  assign out[571] = (in == 10'd571) ? 1'b1 : 1'b0;
  assign out[572] = (in == 10'd572) ? 1'b1 : 1'b0;
  assign out[573] = (in == 10'd573) ? 1'b1 : 1'b0;
  assign out[574] = (in == 10'd574) ? 1'b1 : 1'b0;
  assign out[575] = (in == 10'd575) ? 1'b1 : 1'b0;
  assign out[576] = (in == 10'd576) ? 1'b1 : 1'b0;
  assign out[577] = (in == 10'd577) ? 1'b1 : 1'b0;
  assign out[578] = (in == 10'd578) ? 1'b1 : 1'b0;
  assign out[579] = (in == 10'd579) ? 1'b1 : 1'b0;
  assign out[580] = (in == 10'd580) ? 1'b1 : 1'b0;
  assign out[581] = (in == 10'd581) ? 1'b1 : 1'b0;
  assign out[582] = (in == 10'd582) ? 1'b1 : 1'b0;
  assign out[583] = (in == 10'd583) ? 1'b1 : 1'b0;
  assign out[584] = (in == 10'd584) ? 1'b1 : 1'b0;
  assign out[585] = (in == 10'd585) ? 1'b1 : 1'b0;
  assign out[586] = (in == 10'd586) ? 1'b1 : 1'b0;
  assign out[587] = (in == 10'd587) ? 1'b1 : 1'b0;
  assign out[588] = (in == 10'd588) ? 1'b1 : 1'b0;
  assign out[589] = (in == 10'd589) ? 1'b1 : 1'b0;
  assign out[590] = (in == 10'd590) ? 1'b1 : 1'b0;
  assign out[591] = (in == 10'd591) ? 1'b1 : 1'b0;
  assign out[592] = (in == 10'd592) ? 1'b1 : 1'b0;
  assign out[593] = (in == 10'd593) ? 1'b1 : 1'b0;
  assign out[594] = (in == 10'd594) ? 1'b1 : 1'b0;
  assign out[595] = (in == 10'd595) ? 1'b1 : 1'b0;
  assign out[596] = (in == 10'd596) ? 1'b1 : 1'b0;
  assign out[597] = (in == 10'd597) ? 1'b1 : 1'b0;
  assign out[598] = (in == 10'd598) ? 1'b1 : 1'b0;
  assign out[599] = (in == 10'd599) ? 1'b1 : 1'b0;
  assign out[600] = (in == 10'd600) ? 1'b1 : 1'b0;
  assign out[601] = (in == 10'd601) ? 1'b1 : 1'b0;
  assign out[602] = (in == 10'd602) ? 1'b1 : 1'b0;
  assign out[603] = (in == 10'd603) ? 1'b1 : 1'b0;
  assign out[604] = (in == 10'd604) ? 1'b1 : 1'b0;
  assign out[605] = (in == 10'd605) ? 1'b1 : 1'b0;
  assign out[606] = (in == 10'd606) ? 1'b1 : 1'b0;
  assign out[607] = (in == 10'd607) ? 1'b1 : 1'b0;
  assign out[608] = (in == 10'd608) ? 1'b1 : 1'b0;
  assign out[609] = (in == 10'd609) ? 1'b1 : 1'b0;
  assign out[610] = (in == 10'd610) ? 1'b1 : 1'b0;
  assign out[611] = (in == 10'd611) ? 1'b1 : 1'b0;
  assign out[612] = (in == 10'd612) ? 1'b1 : 1'b0;
  assign out[613] = (in == 10'd613) ? 1'b1 : 1'b0;
  assign out[614] = (in == 10'd614) ? 1'b1 : 1'b0;
  assign out[615] = (in == 10'd615) ? 1'b1 : 1'b0;
  assign out[616] = (in == 10'd616) ? 1'b1 : 1'b0;
  assign out[617] = (in == 10'd617) ? 1'b1 : 1'b0;
  assign out[618] = (in == 10'd618) ? 1'b1 : 1'b0;
  assign out[619] = (in == 10'd619) ? 1'b1 : 1'b0;
  assign out[620] = (in == 10'd620) ? 1'b1 : 1'b0;
  assign out[621] = (in == 10'd621) ? 1'b1 : 1'b0;
  assign out[622] = (in == 10'd622) ? 1'b1 : 1'b0;
  assign out[623] = (in == 10'd623) ? 1'b1 : 1'b0;
  assign out[624] = (in == 10'd624) ? 1'b1 : 1'b0;
  assign out[625] = (in == 10'd625) ? 1'b1 : 1'b0;
  assign out[626] = (in == 10'd626) ? 1'b1 : 1'b0;
  assign out[627] = (in == 10'd627) ? 1'b1 : 1'b0;
  assign out[628] = (in == 10'd628) ? 1'b1 : 1'b0;
  assign out[629] = (in == 10'd629) ? 1'b1 : 1'b0;
  assign out[630] = (in == 10'd630) ? 1'b1 : 1'b0;
  assign out[631] = (in == 10'd631) ? 1'b1 : 1'b0;
  assign out[632] = (in == 10'd632) ? 1'b1 : 1'b0;
  assign out[633] = (in == 10'd633) ? 1'b1 : 1'b0;
  assign out[634] = (in == 10'd634) ? 1'b1 : 1'b0;
  assign out[635] = (in == 10'd635) ? 1'b1 : 1'b0;
  assign out[636] = (in == 10'd636) ? 1'b1 : 1'b0;
  assign out[637] = (in == 10'd637) ? 1'b1 : 1'b0;
  assign out[638] = (in == 10'd638) ? 1'b1 : 1'b0;
  assign out[639] = (in == 10'd639) ? 1'b1 : 1'b0;
  assign out[640] = (in == 10'd640) ? 1'b1 : 1'b0;
  assign out[641] = (in == 10'd641) ? 1'b1 : 1'b0;
  assign out[642] = (in == 10'd642) ? 1'b1 : 1'b0;
  assign out[643] = (in == 10'd643) ? 1'b1 : 1'b0;
  assign out[644] = (in == 10'd644) ? 1'b1 : 1'b0;
  assign out[645] = (in == 10'd645) ? 1'b1 : 1'b0;
  assign out[646] = (in == 10'd646) ? 1'b1 : 1'b0;
  assign out[647] = (in == 10'd647) ? 1'b1 : 1'b0;
  assign out[648] = (in == 10'd648) ? 1'b1 : 1'b0;
  assign out[649] = (in == 10'd649) ? 1'b1 : 1'b0;
  assign out[650] = (in == 10'd650) ? 1'b1 : 1'b0;
  assign out[651] = (in == 10'd651) ? 1'b1 : 1'b0;
  assign out[652] = (in == 10'd652) ? 1'b1 : 1'b0;
  assign out[653] = (in == 10'd653) ? 1'b1 : 1'b0;
  assign out[654] = (in == 10'd654) ? 1'b1 : 1'b0;
  assign out[655] = (in == 10'd655) ? 1'b1 : 1'b0;
  assign out[656] = (in == 10'd656) ? 1'b1 : 1'b0;
  assign out[657] = (in == 10'd657) ? 1'b1 : 1'b0;
  assign out[658] = (in == 10'd658) ? 1'b1 : 1'b0;
  assign out[659] = (in == 10'd659) ? 1'b1 : 1'b0;
  assign out[660] = (in == 10'd660) ? 1'b1 : 1'b0;
  assign out[661] = (in == 10'd661) ? 1'b1 : 1'b0;
  assign out[662] = (in == 10'd662) ? 1'b1 : 1'b0;
  assign out[663] = (in == 10'd663) ? 1'b1 : 1'b0;
  assign out[664] = (in == 10'd664) ? 1'b1 : 1'b0;
  assign out[665] = (in == 10'd665) ? 1'b1 : 1'b0;
  assign out[666] = (in == 10'd666) ? 1'b1 : 1'b0;
  assign out[667] = (in == 10'd667) ? 1'b1 : 1'b0;
  assign out[668] = (in == 10'd668) ? 1'b1 : 1'b0;
  assign out[669] = (in == 10'd669) ? 1'b1 : 1'b0;
  assign out[670] = (in == 10'd670) ? 1'b1 : 1'b0;
  assign out[671] = (in == 10'd671) ? 1'b1 : 1'b0;
  assign out[672] = (in == 10'd672) ? 1'b1 : 1'b0;
  assign out[673] = (in == 10'd673) ? 1'b1 : 1'b0;
  assign out[674] = (in == 10'd674) ? 1'b1 : 1'b0;
  assign out[675] = (in == 10'd675) ? 1'b1 : 1'b0;
  assign out[676] = (in == 10'd676) ? 1'b1 : 1'b0;
  assign out[677] = (in == 10'd677) ? 1'b1 : 1'b0;
  assign out[678] = (in == 10'd678) ? 1'b1 : 1'b0;
  assign out[679] = (in == 10'd679) ? 1'b1 : 1'b0;
  assign out[680] = (in == 10'd680) ? 1'b1 : 1'b0;
  assign out[681] = (in == 10'd681) ? 1'b1 : 1'b0;
  assign out[682] = (in == 10'd682) ? 1'b1 : 1'b0;
  assign out[683] = (in == 10'd683) ? 1'b1 : 1'b0;
  assign out[684] = (in == 10'd684) ? 1'b1 : 1'b0;
  assign out[685] = (in == 10'd685) ? 1'b1 : 1'b0;
  assign out[686] = (in == 10'd686) ? 1'b1 : 1'b0;
  assign out[687] = (in == 10'd687) ? 1'b1 : 1'b0;
  assign out[688] = (in == 10'd688) ? 1'b1 : 1'b0;
  assign out[689] = (in == 10'd689) ? 1'b1 : 1'b0;
  assign out[690] = (in == 10'd690) ? 1'b1 : 1'b0;
  assign out[691] = (in == 10'd691) ? 1'b1 : 1'b0;
  assign out[692] = (in == 10'd692) ? 1'b1 : 1'b0;
  assign out[693] = (in == 10'd693) ? 1'b1 : 1'b0;
  assign out[694] = (in == 10'd694) ? 1'b1 : 1'b0;
  assign out[695] = (in == 10'd695) ? 1'b1 : 1'b0;
  assign out[696] = (in == 10'd696) ? 1'b1 : 1'b0;
  assign out[697] = (in == 10'd697) ? 1'b1 : 1'b0;
  assign out[698] = (in == 10'd698) ? 1'b1 : 1'b0;
  assign out[699] = (in == 10'd699) ? 1'b1 : 1'b0;
  assign out[700] = (in == 10'd700) ? 1'b1 : 1'b0;
  assign out[701] = (in == 10'd701) ? 1'b1 : 1'b0;
  assign out[702] = (in == 10'd702) ? 1'b1 : 1'b0;
  assign out[703] = (in == 10'd703) ? 1'b1 : 1'b0;
  assign out[704] = (in == 10'd704) ? 1'b1 : 1'b0;
  assign out[705] = (in == 10'd705) ? 1'b1 : 1'b0;
  assign out[706] = (in == 10'd706) ? 1'b1 : 1'b0;
  assign out[707] = (in == 10'd707) ? 1'b1 : 1'b0;
  assign out[708] = (in == 10'd708) ? 1'b1 : 1'b0;
  assign out[709] = (in == 10'd709) ? 1'b1 : 1'b0;
  assign out[710] = (in == 10'd710) ? 1'b1 : 1'b0;
  assign out[711] = (in == 10'd711) ? 1'b1 : 1'b0;
  assign out[712] = (in == 10'd712) ? 1'b1 : 1'b0;
  assign out[713] = (in == 10'd713) ? 1'b1 : 1'b0;
  assign out[714] = (in == 10'd714) ? 1'b1 : 1'b0;
  assign out[715] = (in == 10'd715) ? 1'b1 : 1'b0;
  assign out[716] = (in == 10'd716) ? 1'b1 : 1'b0;
  assign out[717] = (in == 10'd717) ? 1'b1 : 1'b0;
  assign out[718] = (in == 10'd718) ? 1'b1 : 1'b0;
  assign out[719] = (in == 10'd719) ? 1'b1 : 1'b0;
  assign out[720] = (in == 10'd720) ? 1'b1 : 1'b0;
  assign out[721] = (in == 10'd721) ? 1'b1 : 1'b0;
  assign out[722] = (in == 10'd722) ? 1'b1 : 1'b0;
  assign out[723] = (in == 10'd723) ? 1'b1 : 1'b0;
  assign out[724] = (in == 10'd724) ? 1'b1 : 1'b0;
  assign out[725] = (in == 10'd725) ? 1'b1 : 1'b0;
  assign out[726] = (in == 10'd726) ? 1'b1 : 1'b0;
  assign out[727] = (in == 10'd727) ? 1'b1 : 1'b0;
  assign out[728] = (in == 10'd728) ? 1'b1 : 1'b0;
  assign out[729] = (in == 10'd729) ? 1'b1 : 1'b0;
  assign out[730] = (in == 10'd730) ? 1'b1 : 1'b0;
  assign out[731] = (in == 10'd731) ? 1'b1 : 1'b0;
  assign out[732] = (in == 10'd732) ? 1'b1 : 1'b0;
  assign out[733] = (in == 10'd733) ? 1'b1 : 1'b0;
  assign out[734] = (in == 10'd734) ? 1'b1 : 1'b0;
  assign out[735] = (in == 10'd735) ? 1'b1 : 1'b0;
  assign out[736] = (in == 10'd736) ? 1'b1 : 1'b0;
  assign out[737] = (in == 10'd737) ? 1'b1 : 1'b0;
  assign out[738] = (in == 10'd738) ? 1'b1 : 1'b0;
  assign out[739] = (in == 10'd739) ? 1'b1 : 1'b0;
  assign out[740] = (in == 10'd740) ? 1'b1 : 1'b0;
  assign out[741] = (in == 10'd741) ? 1'b1 : 1'b0;
  assign out[742] = (in == 10'd742) ? 1'b1 : 1'b0;
  assign out[743] = (in == 10'd743) ? 1'b1 : 1'b0;
  assign out[744] = (in == 10'd744) ? 1'b1 : 1'b0;
  assign out[745] = (in == 10'd745) ? 1'b1 : 1'b0;
  assign out[746] = (in == 10'd746) ? 1'b1 : 1'b0;
  assign out[747] = (in == 10'd747) ? 1'b1 : 1'b0;
  assign out[748] = (in == 10'd748) ? 1'b1 : 1'b0;
  assign out[749] = (in == 10'd749) ? 1'b1 : 1'b0;
  assign out[750] = (in == 10'd750) ? 1'b1 : 1'b0;
  assign out[751] = (in == 10'd751) ? 1'b1 : 1'b0;
  assign out[752] = (in == 10'd752) ? 1'b1 : 1'b0;
  assign out[753] = (in == 10'd753) ? 1'b1 : 1'b0;
  assign out[754] = (in == 10'd754) ? 1'b1 : 1'b0;
  assign out[755] = (in == 10'd755) ? 1'b1 : 1'b0;
  assign out[756] = (in == 10'd756) ? 1'b1 : 1'b0;
  assign out[757] = (in == 10'd757) ? 1'b1 : 1'b0;
  assign out[758] = (in == 10'd758) ? 1'b1 : 1'b0;
  assign out[759] = (in == 10'd759) ? 1'b1 : 1'b0;
  assign out[760] = (in == 10'd760) ? 1'b1 : 1'b0;
  assign out[761] = (in == 10'd761) ? 1'b1 : 1'b0;
  assign out[762] = (in == 10'd762) ? 1'b1 : 1'b0;
  assign out[763] = (in == 10'd763) ? 1'b1 : 1'b0;
  assign out[764] = (in == 10'd764) ? 1'b1 : 1'b0;
  assign out[765] = (in == 10'd765) ? 1'b1 : 1'b0;
  assign out[766] = (in == 10'd766) ? 1'b1 : 1'b0;
  assign out[767] = (in == 10'd767) ? 1'b1 : 1'b0;
  assign out[768] = (in == 10'd768) ? 1'b1 : 1'b0;
  assign out[769] = (in == 10'd769) ? 1'b1 : 1'b0;
  assign out[770] = (in == 10'd770) ? 1'b1 : 1'b0;
  assign out[771] = (in == 10'd771) ? 1'b1 : 1'b0;
  assign out[772] = (in == 10'd772) ? 1'b1 : 1'b0;
  assign out[773] = (in == 10'd773) ? 1'b1 : 1'b0;
  assign out[774] = (in == 10'd774) ? 1'b1 : 1'b0;
  assign out[775] = (in == 10'd775) ? 1'b1 : 1'b0;
  assign out[776] = (in == 10'd776) ? 1'b1 : 1'b0;
  assign out[777] = (in == 10'd777) ? 1'b1 : 1'b0;
  assign out[778] = (in == 10'd778) ? 1'b1 : 1'b0;
  assign out[779] = (in == 10'd779) ? 1'b1 : 1'b0;
  assign out[780] = (in == 10'd780) ? 1'b1 : 1'b0;
  assign out[781] = (in == 10'd781) ? 1'b1 : 1'b0;
  assign out[782] = (in == 10'd782) ? 1'b1 : 1'b0;
  assign out[783] = (in == 10'd783) ? 1'b1 : 1'b0;
  assign out[784] = (in == 10'd784) ? 1'b1 : 1'b0;
  assign out[785] = (in == 10'd785) ? 1'b1 : 1'b0;
  assign out[786] = (in == 10'd786) ? 1'b1 : 1'b0;
  assign out[787] = (in == 10'd787) ? 1'b1 : 1'b0;
  assign out[788] = (in == 10'd788) ? 1'b1 : 1'b0;
  assign out[789] = (in == 10'd789) ? 1'b1 : 1'b0;
  assign out[790] = (in == 10'd790) ? 1'b1 : 1'b0;
  assign out[791] = (in == 10'd791) ? 1'b1 : 1'b0;
  assign out[792] = (in == 10'd792) ? 1'b1 : 1'b0;
  assign out[793] = (in == 10'd793) ? 1'b1 : 1'b0;
  assign out[794] = (in == 10'd794) ? 1'b1 : 1'b0;
  assign out[795] = (in == 10'd795) ? 1'b1 : 1'b0;
  assign out[796] = (in == 10'd796) ? 1'b1 : 1'b0;
  assign out[797] = (in == 10'd797) ? 1'b1 : 1'b0;
  assign out[798] = (in == 10'd798) ? 1'b1 : 1'b0;
  assign out[799] = (in == 10'd799) ? 1'b1 : 1'b0;
  assign out[800] = (in == 10'd800) ? 1'b1 : 1'b0;
  assign out[801] = (in == 10'd801) ? 1'b1 : 1'b0;
  assign out[802] = (in == 10'd802) ? 1'b1 : 1'b0;
  assign out[803] = (in == 10'd803) ? 1'b1 : 1'b0;
  assign out[804] = (in == 10'd804) ? 1'b1 : 1'b0;
  assign out[805] = (in == 10'd805) ? 1'b1 : 1'b0;
  assign out[806] = (in == 10'd806) ? 1'b1 : 1'b0;
  assign out[807] = (in == 10'd807) ? 1'b1 : 1'b0;
  assign out[808] = (in == 10'd808) ? 1'b1 : 1'b0;
  assign out[809] = (in == 10'd809) ? 1'b1 : 1'b0;
  assign out[810] = (in == 10'd810) ? 1'b1 : 1'b0;
  assign out[811] = (in == 10'd811) ? 1'b1 : 1'b0;
  assign out[812] = (in == 10'd812) ? 1'b1 : 1'b0;
  assign out[813] = (in == 10'd813) ? 1'b1 : 1'b0;
  assign out[814] = (in == 10'd814) ? 1'b1 : 1'b0;
  assign out[815] = (in == 10'd815) ? 1'b1 : 1'b0;
  assign out[816] = (in == 10'd816) ? 1'b1 : 1'b0;
  assign out[817] = (in == 10'd817) ? 1'b1 : 1'b0;
  assign out[818] = (in == 10'd818) ? 1'b1 : 1'b0;
  assign out[819] = (in == 10'd819) ? 1'b1 : 1'b0;
  assign out[820] = (in == 10'd820) ? 1'b1 : 1'b0;
  assign out[821] = (in == 10'd821) ? 1'b1 : 1'b0;
  assign out[822] = (in == 10'd822) ? 1'b1 : 1'b0;
  assign out[823] = (in == 10'd823) ? 1'b1 : 1'b0;
  assign out[824] = (in == 10'd824) ? 1'b1 : 1'b0;
  assign out[825] = (in == 10'd825) ? 1'b1 : 1'b0;
  assign out[826] = (in == 10'd826) ? 1'b1 : 1'b0;
  assign out[827] = (in == 10'd827) ? 1'b1 : 1'b0;
  assign out[828] = (in == 10'd828) ? 1'b1 : 1'b0;
  assign out[829] = (in == 10'd829) ? 1'b1 : 1'b0;
  assign out[830] = (in == 10'd830) ? 1'b1 : 1'b0;
  assign out[831] = (in == 10'd831) ? 1'b1 : 1'b0;
  assign out[832] = (in == 10'd832) ? 1'b1 : 1'b0;
  assign out[833] = (in == 10'd833) ? 1'b1 : 1'b0;
  assign out[834] = (in == 10'd834) ? 1'b1 : 1'b0;
  assign out[835] = (in == 10'd835) ? 1'b1 : 1'b0;
  assign out[836] = (in == 10'd836) ? 1'b1 : 1'b0;
  assign out[837] = (in == 10'd837) ? 1'b1 : 1'b0;
  assign out[838] = (in == 10'd838) ? 1'b1 : 1'b0;
  assign out[839] = (in == 10'd839) ? 1'b1 : 1'b0;
  assign out[840] = (in == 10'd840) ? 1'b1 : 1'b0;
  assign out[841] = (in == 10'd841) ? 1'b1 : 1'b0;
  assign out[842] = (in == 10'd842) ? 1'b1 : 1'b0;
  assign out[843] = (in == 10'd843) ? 1'b1 : 1'b0;
  assign out[844] = (in == 10'd844) ? 1'b1 : 1'b0;
  assign out[845] = (in == 10'd845) ? 1'b1 : 1'b0;
  assign out[846] = (in == 10'd846) ? 1'b1 : 1'b0;
  assign out[847] = (in == 10'd847) ? 1'b1 : 1'b0;
  assign out[848] = (in == 10'd848) ? 1'b1 : 1'b0;
  assign out[849] = (in == 10'd849) ? 1'b1 : 1'b0;
  assign out[850] = (in == 10'd850) ? 1'b1 : 1'b0;
  assign out[851] = (in == 10'd851) ? 1'b1 : 1'b0;
  assign out[852] = (in == 10'd852) ? 1'b1 : 1'b0;
  assign out[853] = (in == 10'd853) ? 1'b1 : 1'b0;
  assign out[854] = (in == 10'd854) ? 1'b1 : 1'b0;
  assign out[855] = (in == 10'd855) ? 1'b1 : 1'b0;
  assign out[856] = (in == 10'd856) ? 1'b1 : 1'b0;
  assign out[857] = (in == 10'd857) ? 1'b1 : 1'b0;
  assign out[858] = (in == 10'd858) ? 1'b1 : 1'b0;
  assign out[859] = (in == 10'd859) ? 1'b1 : 1'b0;
  assign out[860] = (in == 10'd860) ? 1'b1 : 1'b0;
  assign out[861] = (in == 10'd861) ? 1'b1 : 1'b0;
  assign out[862] = (in == 10'd862) ? 1'b1 : 1'b0;
  assign out[863] = (in == 10'd863) ? 1'b1 : 1'b0;
  assign out[864] = (in == 10'd864) ? 1'b1 : 1'b0;
  assign out[865] = (in == 10'd865) ? 1'b1 : 1'b0;
  assign out[866] = (in == 10'd866) ? 1'b1 : 1'b0;
  assign out[867] = (in == 10'd867) ? 1'b1 : 1'b0;
  assign out[868] = (in == 10'd868) ? 1'b1 : 1'b0;
  assign out[869] = (in == 10'd869) ? 1'b1 : 1'b0;
  assign out[870] = (in == 10'd870) ? 1'b1 : 1'b0;
  assign out[871] = (in == 10'd871) ? 1'b1 : 1'b0;
  assign out[872] = (in == 10'd872) ? 1'b1 : 1'b0;
  assign out[873] = (in == 10'd873) ? 1'b1 : 1'b0;
  assign out[874] = (in == 10'd874) ? 1'b1 : 1'b0;
  assign out[875] = (in == 10'd875) ? 1'b1 : 1'b0;
  assign out[876] = (in == 10'd876) ? 1'b1 : 1'b0;
  assign out[877] = (in == 10'd877) ? 1'b1 : 1'b0;
  assign out[878] = (in == 10'd878) ? 1'b1 : 1'b0;
  assign out[879] = (in == 10'd879) ? 1'b1 : 1'b0;
  assign out[880] = (in == 10'd880) ? 1'b1 : 1'b0;
  assign out[881] = (in == 10'd881) ? 1'b1 : 1'b0;
  assign out[882] = (in == 10'd882) ? 1'b1 : 1'b0;
  assign out[883] = (in == 10'd883) ? 1'b1 : 1'b0;
  assign out[884] = (in == 10'd884) ? 1'b1 : 1'b0;
  assign out[885] = (in == 10'd885) ? 1'b1 : 1'b0;
  assign out[886] = (in == 10'd886) ? 1'b1 : 1'b0;
  assign out[887] = (in == 10'd887) ? 1'b1 : 1'b0;
  assign out[888] = (in == 10'd888) ? 1'b1 : 1'b0;
  assign out[889] = (in == 10'd889) ? 1'b1 : 1'b0;
  assign out[890] = (in == 10'd890) ? 1'b1 : 1'b0;
  assign out[891] = (in == 10'd891) ? 1'b1 : 1'b0;
  assign out[892] = (in == 10'd892) ? 1'b1 : 1'b0;
  assign out[893] = (in == 10'd893) ? 1'b1 : 1'b0;
  assign out[894] = (in == 10'd894) ? 1'b1 : 1'b0;
  assign out[895] = (in == 10'd895) ? 1'b1 : 1'b0;
  assign out[896] = (in == 10'd896) ? 1'b1 : 1'b0;
  assign out[897] = (in == 10'd897) ? 1'b1 : 1'b0;
  assign out[898] = (in == 10'd898) ? 1'b1 : 1'b0;
  assign out[899] = (in == 10'd899) ? 1'b1 : 1'b0;
  assign out[900] = (in == 10'd900) ? 1'b1 : 1'b0;
  assign out[901] = (in == 10'd901) ? 1'b1 : 1'b0;
  assign out[902] = (in == 10'd902) ? 1'b1 : 1'b0;
  assign out[903] = (in == 10'd903) ? 1'b1 : 1'b0;
  assign out[904] = (in == 10'd904) ? 1'b1 : 1'b0;
  assign out[905] = (in == 10'd905) ? 1'b1 : 1'b0;
  assign out[906] = (in == 10'd906) ? 1'b1 : 1'b0;
  assign out[907] = (in == 10'd907) ? 1'b1 : 1'b0;
  assign out[908] = (in == 10'd908) ? 1'b1 : 1'b0;
  assign out[909] = (in == 10'd909) ? 1'b1 : 1'b0;
  assign out[910] = (in == 10'd910) ? 1'b1 : 1'b0;
  assign out[911] = (in == 10'd911) ? 1'b1 : 1'b0;
  assign out[912] = (in == 10'd912) ? 1'b1 : 1'b0;
  assign out[913] = (in == 10'd913) ? 1'b1 : 1'b0;
  assign out[914] = (in == 10'd914) ? 1'b1 : 1'b0;
  assign out[915] = (in == 10'd915) ? 1'b1 : 1'b0;
  assign out[916] = (in == 10'd916) ? 1'b1 : 1'b0;
  assign out[917] = (in == 10'd917) ? 1'b1 : 1'b0;
  assign out[918] = (in == 10'd918) ? 1'b1 : 1'b0;
  assign out[919] = (in == 10'd919) ? 1'b1 : 1'b0;
  assign out[920] = (in == 10'd920) ? 1'b1 : 1'b0;
  assign out[921] = (in == 10'd921) ? 1'b1 : 1'b0;
  assign out[922] = (in == 10'd922) ? 1'b1 : 1'b0;
  assign out[923] = (in == 10'd923) ? 1'b1 : 1'b0;
  assign out[924] = (in == 10'd924) ? 1'b1 : 1'b0;
  assign out[925] = (in == 10'd925) ? 1'b1 : 1'b0;
  assign out[926] = (in == 10'd926) ? 1'b1 : 1'b0;
  assign out[927] = (in == 10'd927) ? 1'b1 : 1'b0;
  assign out[928] = (in == 10'd928) ? 1'b1 : 1'b0;
  assign out[929] = (in == 10'd929) ? 1'b1 : 1'b0;
  assign out[930] = (in == 10'd930) ? 1'b1 : 1'b0;
  assign out[931] = (in == 10'd931) ? 1'b1 : 1'b0;
  assign out[932] = (in == 10'd932) ? 1'b1 : 1'b0;
  assign out[933] = (in == 10'd933) ? 1'b1 : 1'b0;
  assign out[934] = (in == 10'd934) ? 1'b1 : 1'b0;
  assign out[935] = (in == 10'd935) ? 1'b1 : 1'b0;
  assign out[936] = (in == 10'd936) ? 1'b1 : 1'b0;
  assign out[937] = (in == 10'd937) ? 1'b1 : 1'b0;
  assign out[938] = (in == 10'd938) ? 1'b1 : 1'b0;
  assign out[939] = (in == 10'd939) ? 1'b1 : 1'b0;
  assign out[940] = (in == 10'd940) ? 1'b1 : 1'b0;
  assign out[941] = (in == 10'd941) ? 1'b1 : 1'b0;
  assign out[942] = (in == 10'd942) ? 1'b1 : 1'b0;
  assign out[943] = (in == 10'd943) ? 1'b1 : 1'b0;
  assign out[944] = (in == 10'd944) ? 1'b1 : 1'b0;
  assign out[945] = (in == 10'd945) ? 1'b1 : 1'b0;
  assign out[946] = (in == 10'd946) ? 1'b1 : 1'b0;
  assign out[947] = (in == 10'd947) ? 1'b1 : 1'b0;
  assign out[948] = (in == 10'd948) ? 1'b1 : 1'b0;
  assign out[949] = (in == 10'd949) ? 1'b1 : 1'b0;
  assign out[950] = (in == 10'd950) ? 1'b1 : 1'b0;
  assign out[951] = (in == 10'd951) ? 1'b1 : 1'b0;
  assign out[952] = (in == 10'd952) ? 1'b1 : 1'b0;
  assign out[953] = (in == 10'd953) ? 1'b1 : 1'b0;
  assign out[954] = (in == 10'd954) ? 1'b1 : 1'b0;
  assign out[955] = (in == 10'd955) ? 1'b1 : 1'b0;
  assign out[956] = (in == 10'd956) ? 1'b1 : 1'b0;
  assign out[957] = (in == 10'd957) ? 1'b1 : 1'b0;
  assign out[958] = (in == 10'd958) ? 1'b1 : 1'b0;
  assign out[959] = (in == 10'd959) ? 1'b1 : 1'b0;
  assign out[960] = (in == 10'd960) ? 1'b1 : 1'b0;
  assign out[961] = (in == 10'd961) ? 1'b1 : 1'b0;
  assign out[962] = (in == 10'd962) ? 1'b1 : 1'b0;
  assign out[963] = (in == 10'd963) ? 1'b1 : 1'b0;
  assign out[964] = (in == 10'd964) ? 1'b1 : 1'b0;
  assign out[965] = (in == 10'd965) ? 1'b1 : 1'b0;
  assign out[966] = (in == 10'd966) ? 1'b1 : 1'b0;
  assign out[967] = (in == 10'd967) ? 1'b1 : 1'b0;
  assign out[968] = (in == 10'd968) ? 1'b1 : 1'b0;
  assign out[969] = (in == 10'd969) ? 1'b1 : 1'b0;
  assign out[970] = (in == 10'd970) ? 1'b1 : 1'b0;
  assign out[971] = (in == 10'd971) ? 1'b1 : 1'b0;
  assign out[972] = (in == 10'd972) ? 1'b1 : 1'b0;
  assign out[973] = (in == 10'd973) ? 1'b1 : 1'b0;
  assign out[974] = (in == 10'd974) ? 1'b1 : 1'b0;
  assign out[975] = (in == 10'd975) ? 1'b1 : 1'b0;
  assign out[976] = (in == 10'd976) ? 1'b1 : 1'b0;
  assign out[977] = (in == 10'd977) ? 1'b1 : 1'b0;
  assign out[978] = (in == 10'd978) ? 1'b1 : 1'b0;
  assign out[979] = (in == 10'd979) ? 1'b1 : 1'b0;
  assign out[980] = (in == 10'd980) ? 1'b1 : 1'b0;
  assign out[981] = (in == 10'd981) ? 1'b1 : 1'b0;
  assign out[982] = (in == 10'd982) ? 1'b1 : 1'b0;
  assign out[983] = (in == 10'd983) ? 1'b1 : 1'b0;
  assign out[984] = (in == 10'd984) ? 1'b1 : 1'b0;
  assign out[985] = (in == 10'd985) ? 1'b1 : 1'b0;
  assign out[986] = (in == 10'd986) ? 1'b1 : 1'b0;
  assign out[987] = (in == 10'd987) ? 1'b1 : 1'b0;
  assign out[988] = (in == 10'd988) ? 1'b1 : 1'b0;
  assign out[989] = (in == 10'd989) ? 1'b1 : 1'b0;
  assign out[990] = (in == 10'd990) ? 1'b1 : 1'b0;
  assign out[991] = (in == 10'd991) ? 1'b1 : 1'b0;
  assign out[992] = (in == 10'd992) ? 1'b1 : 1'b0;
  assign out[993] = (in == 10'd993) ? 1'b1 : 1'b0;
  assign out[994] = (in == 10'd994) ? 1'b1 : 1'b0;
  assign out[995] = (in == 10'd995) ? 1'b1 : 1'b0;
  assign out[996] = (in == 10'd996) ? 1'b1 : 1'b0;
  assign out[997] = (in == 10'd997) ? 1'b1 : 1'b0;
  assign out[998] = (in == 10'd998) ? 1'b1 : 1'b0;
  assign out[999] = (in == 10'd999) ? 1'b1 : 1'b0;
  assign out[1000] = (in == 10'd1000) ? 1'b1 : 1'b0;
  assign out[1001] = (in == 10'd1001) ? 1'b1 : 1'b0;
  assign out[1002] = (in == 10'd1002) ? 1'b1 : 1'b0;
  assign out[1003] = (in == 10'd1003) ? 1'b1 : 1'b0;
  assign out[1004] = (in == 10'd1004) ? 1'b1 : 1'b0;
  assign out[1005] = (in == 10'd1005) ? 1'b1 : 1'b0;
  assign out[1006] = (in == 10'd1006) ? 1'b1 : 1'b0;
  assign out[1007] = (in == 10'd1007) ? 1'b1 : 1'b0;
  assign out[1008] = (in == 10'd1008) ? 1'b1 : 1'b0;
  assign out[1009] = (in == 10'd1009) ? 1'b1 : 1'b0;
  assign out[1010] = (in == 10'd1010) ? 1'b1 : 1'b0;
  assign out[1011] = (in == 10'd1011) ? 1'b1 : 1'b0;
  assign out[1012] = (in == 10'd1012) ? 1'b1 : 1'b0;
  assign out[1013] = (in == 10'd1013) ? 1'b1 : 1'b0;
  assign out[1014] = (in == 10'd1014) ? 1'b1 : 1'b0;
  assign out[1015] = (in == 10'd1015) ? 1'b1 : 1'b0;
  assign out[1016] = (in == 10'd1016) ? 1'b1 : 1'b0;
  assign out[1017] = (in == 10'd1017) ? 1'b1 : 1'b0;
  assign out[1018] = (in == 10'd1018) ? 1'b1 : 1'b0;
  assign out[1019] = (in == 10'd1019) ? 1'b1 : 1'b0;
  assign out[1020] = (in == 10'd1020) ? 1'b1 : 1'b0;
  assign out[1021] = (in == 10'd1021) ? 1'b1 : 1'b0;
  assign out[1022] = (in == 10'd1022) ? 1'b1 : 1'b0;
  assign out[1023] = (in == 10'd1023) ? 1'b1 : 1'b0;
endmodule
