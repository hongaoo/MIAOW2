`define FPGA_BUILD 1
`include "alu_definitions.v"
`include "decode_definitions.v"
`include "issue_definitions.v"
`include "lsu_definitions.v"
`include "global_definitions.v"
module reg_128x32b_3r_3w
(
  rd0_data, rd1_data, rd2_data,
  clk,
  rd0_addr, rd1_addr, rd2_addr,
  wr0_addr, wr1_addr, wr2_addr,
  wr0_en, wr1_en, wr2_en, wr0_data, wr1_data, wr2_data
);
input clk;

output [31:0] rd0_data;
output [31:0] rd1_data;
output [31:0] rd2_data;

input [6:0] rd0_addr;
input [6:0] rd1_addr;
input [6:0] rd2_addr;

input [6:0] wr0_addr;
input [6:0] wr1_addr;
input [6:0] wr2_addr;

input wr0_en;
input wr1_en;
input wr2_en;

input [31:0] wr0_data;
input [31:0] wr1_data;
input [31:0] wr2_data;

wire [4095:0] word_out;
wire [4095:0] word_in;
wire [127:0] wr_en_word;

wire [127:0] wr0_word_select;
wire [127:0] wr1_word_select;
wire [127:0] wr2_word_select;
wire [127:0] wr0_word_enable;
wire [127:0] wr1_word_enable;
wire [127:0] wr2_word_enable;

//Register file
flop_32b word[127:0](.out(word_out), .in(word_in), .wr_en(wr_en_word), .clk(clk));

//Muxes for read ports
mux_128x32b_to_1x32b mux_rd_port_0 (.out(rd0_data), .in(word_out), .select(rd0_addr));
mux_128x32b_to_1x32b mux_rd_port_1 (.out(rd1_data), .in(word_out), .select(rd1_addr));
mux_128x32b_to_1x32b mux_rd_port_2 (.out(rd2_data), .in(word_out), .select(rd2_addr));

//Write port logic
decoder_param #(7,128) decoder_wr_port_0 (.out(wr0_word_select), .in(wr0_addr));
decoder_param #(7,128) decoder_wr_port_1 (.out(wr1_word_select), .in(wr1_addr));
decoder_param #(7,128) decoder_wr_port_2 (.out(wr2_word_select), .in(wr2_addr));
assign wr0_word_enable = {128{wr0_en}} & wr0_word_select;
assign wr1_word_enable = {128{wr1_en}} & wr1_word_select;
assign wr2_word_enable = {128{wr2_en}} & wr2_word_select;
assign wr_en_word = wr0_word_enable | wr1_word_enable | wr2_word_enable;

// %%start_veriperl
// my $i;
// my $low_index;
// my $high_index;
// for($i=0; $i<128; $i=$i+1)
// {
//   $low_index = 32*$i;
//   $high_index = 32*$i+31;
//   print "assign word_in[$high_index:$low_index] = ({wr2_word_enable[$i],wr1_word_enable[$i],wr0_word_enable[$i]} == 3'b001) ? wr0_data : (({wr2_word_enable[$i],wr1_word_enable[$i],wr0_word_enable[$i]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[$i],wr1_word_enable[$i],wr0_word_enable[$i]} == 3'b100)? wr2_data : {32{1'bx}}));\n";
// }
// %%stop_veriperl
assign word_in[31:0] = ({wr2_word_enable[0],wr1_word_enable[0],wr0_word_enable[0]} == 3'b001) ? wr0_data : (({wr2_word_enable[0],wr1_word_enable[0],wr0_word_enable[0]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[0],wr1_word_enable[0],wr0_word_enable[0]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[63:32] = ({wr2_word_enable[1],wr1_word_enable[1],wr0_word_enable[1]} == 3'b001) ? wr0_data : (({wr2_word_enable[1],wr1_word_enable[1],wr0_word_enable[1]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[1],wr1_word_enable[1],wr0_word_enable[1]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[95:64] = ({wr2_word_enable[2],wr1_word_enable[2],wr0_word_enable[2]} == 3'b001) ? wr0_data : (({wr2_word_enable[2],wr1_word_enable[2],wr0_word_enable[2]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[2],wr1_word_enable[2],wr0_word_enable[2]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[127:96] = ({wr2_word_enable[3],wr1_word_enable[3],wr0_word_enable[3]} == 3'b001) ? wr0_data : (({wr2_word_enable[3],wr1_word_enable[3],wr0_word_enable[3]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[3],wr1_word_enable[3],wr0_word_enable[3]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[159:128] = ({wr2_word_enable[4],wr1_word_enable[4],wr0_word_enable[4]} == 3'b001) ? wr0_data : (({wr2_word_enable[4],wr1_word_enable[4],wr0_word_enable[4]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[4],wr1_word_enable[4],wr0_word_enable[4]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[191:160] = ({wr2_word_enable[5],wr1_word_enable[5],wr0_word_enable[5]} == 3'b001) ? wr0_data : (({wr2_word_enable[5],wr1_word_enable[5],wr0_word_enable[5]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[5],wr1_word_enable[5],wr0_word_enable[5]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[223:192] = ({wr2_word_enable[6],wr1_word_enable[6],wr0_word_enable[6]} == 3'b001) ? wr0_data : (({wr2_word_enable[6],wr1_word_enable[6],wr0_word_enable[6]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[6],wr1_word_enable[6],wr0_word_enable[6]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[255:224] = ({wr2_word_enable[7],wr1_word_enable[7],wr0_word_enable[7]} == 3'b001) ? wr0_data : (({wr2_word_enable[7],wr1_word_enable[7],wr0_word_enable[7]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[7],wr1_word_enable[7],wr0_word_enable[7]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[287:256] = ({wr2_word_enable[8],wr1_word_enable[8],wr0_word_enable[8]} == 3'b001) ? wr0_data : (({wr2_word_enable[8],wr1_word_enable[8],wr0_word_enable[8]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[8],wr1_word_enable[8],wr0_word_enable[8]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[319:288] = ({wr2_word_enable[9],wr1_word_enable[9],wr0_word_enable[9]} == 3'b001) ? wr0_data : (({wr2_word_enable[9],wr1_word_enable[9],wr0_word_enable[9]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[9],wr1_word_enable[9],wr0_word_enable[9]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[351:320] = ({wr2_word_enable[10],wr1_word_enable[10],wr0_word_enable[10]} == 3'b001) ? wr0_data : (({wr2_word_enable[10],wr1_word_enable[10],wr0_word_enable[10]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[10],wr1_word_enable[10],wr0_word_enable[10]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[383:352] = ({wr2_word_enable[11],wr1_word_enable[11],wr0_word_enable[11]} == 3'b001) ? wr0_data : (({wr2_word_enable[11],wr1_word_enable[11],wr0_word_enable[11]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[11],wr1_word_enable[11],wr0_word_enable[11]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[415:384] = ({wr2_word_enable[12],wr1_word_enable[12],wr0_word_enable[12]} == 3'b001) ? wr0_data : (({wr2_word_enable[12],wr1_word_enable[12],wr0_word_enable[12]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[12],wr1_word_enable[12],wr0_word_enable[12]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[447:416] = ({wr2_word_enable[13],wr1_word_enable[13],wr0_word_enable[13]} == 3'b001) ? wr0_data : (({wr2_word_enable[13],wr1_word_enable[13],wr0_word_enable[13]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[13],wr1_word_enable[13],wr0_word_enable[13]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[479:448] = ({wr2_word_enable[14],wr1_word_enable[14],wr0_word_enable[14]} == 3'b001) ? wr0_data : (({wr2_word_enable[14],wr1_word_enable[14],wr0_word_enable[14]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[14],wr1_word_enable[14],wr0_word_enable[14]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[511:480] = ({wr2_word_enable[15],wr1_word_enable[15],wr0_word_enable[15]} == 3'b001) ? wr0_data : (({wr2_word_enable[15],wr1_word_enable[15],wr0_word_enable[15]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[15],wr1_word_enable[15],wr0_word_enable[15]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[543:512] = ({wr2_word_enable[16],wr1_word_enable[16],wr0_word_enable[16]} == 3'b001) ? wr0_data : (({wr2_word_enable[16],wr1_word_enable[16],wr0_word_enable[16]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[16],wr1_word_enable[16],wr0_word_enable[16]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[575:544] = ({wr2_word_enable[17],wr1_word_enable[17],wr0_word_enable[17]} == 3'b001) ? wr0_data : (({wr2_word_enable[17],wr1_word_enable[17],wr0_word_enable[17]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[17],wr1_word_enable[17],wr0_word_enable[17]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[607:576] = ({wr2_word_enable[18],wr1_word_enable[18],wr0_word_enable[18]} == 3'b001) ? wr0_data : (({wr2_word_enable[18],wr1_word_enable[18],wr0_word_enable[18]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[18],wr1_word_enable[18],wr0_word_enable[18]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[639:608] = ({wr2_word_enable[19],wr1_word_enable[19],wr0_word_enable[19]} == 3'b001) ? wr0_data : (({wr2_word_enable[19],wr1_word_enable[19],wr0_word_enable[19]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[19],wr1_word_enable[19],wr0_word_enable[19]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[671:640] = ({wr2_word_enable[20],wr1_word_enable[20],wr0_word_enable[20]} == 3'b001) ? wr0_data : (({wr2_word_enable[20],wr1_word_enable[20],wr0_word_enable[20]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[20],wr1_word_enable[20],wr0_word_enable[20]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[703:672] = ({wr2_word_enable[21],wr1_word_enable[21],wr0_word_enable[21]} == 3'b001) ? wr0_data : (({wr2_word_enable[21],wr1_word_enable[21],wr0_word_enable[21]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[21],wr1_word_enable[21],wr0_word_enable[21]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[735:704] = ({wr2_word_enable[22],wr1_word_enable[22],wr0_word_enable[22]} == 3'b001) ? wr0_data : (({wr2_word_enable[22],wr1_word_enable[22],wr0_word_enable[22]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[22],wr1_word_enable[22],wr0_word_enable[22]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[767:736] = ({wr2_word_enable[23],wr1_word_enable[23],wr0_word_enable[23]} == 3'b001) ? wr0_data : (({wr2_word_enable[23],wr1_word_enable[23],wr0_word_enable[23]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[23],wr1_word_enable[23],wr0_word_enable[23]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[799:768] = ({wr2_word_enable[24],wr1_word_enable[24],wr0_word_enable[24]} == 3'b001) ? wr0_data : (({wr2_word_enable[24],wr1_word_enable[24],wr0_word_enable[24]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[24],wr1_word_enable[24],wr0_word_enable[24]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[831:800] = ({wr2_word_enable[25],wr1_word_enable[25],wr0_word_enable[25]} == 3'b001) ? wr0_data : (({wr2_word_enable[25],wr1_word_enable[25],wr0_word_enable[25]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[25],wr1_word_enable[25],wr0_word_enable[25]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[863:832] = ({wr2_word_enable[26],wr1_word_enable[26],wr0_word_enable[26]} == 3'b001) ? wr0_data : (({wr2_word_enable[26],wr1_word_enable[26],wr0_word_enable[26]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[26],wr1_word_enable[26],wr0_word_enable[26]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[895:864] = ({wr2_word_enable[27],wr1_word_enable[27],wr0_word_enable[27]} == 3'b001) ? wr0_data : (({wr2_word_enable[27],wr1_word_enable[27],wr0_word_enable[27]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[27],wr1_word_enable[27],wr0_word_enable[27]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[927:896] = ({wr2_word_enable[28],wr1_word_enable[28],wr0_word_enable[28]} == 3'b001) ? wr0_data : (({wr2_word_enable[28],wr1_word_enable[28],wr0_word_enable[28]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[28],wr1_word_enable[28],wr0_word_enable[28]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[959:928] = ({wr2_word_enable[29],wr1_word_enable[29],wr0_word_enable[29]} == 3'b001) ? wr0_data : (({wr2_word_enable[29],wr1_word_enable[29],wr0_word_enable[29]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[29],wr1_word_enable[29],wr0_word_enable[29]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[991:960] = ({wr2_word_enable[30],wr1_word_enable[30],wr0_word_enable[30]} == 3'b001) ? wr0_data : (({wr2_word_enable[30],wr1_word_enable[30],wr0_word_enable[30]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[30],wr1_word_enable[30],wr0_word_enable[30]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1023:992] = ({wr2_word_enable[31],wr1_word_enable[31],wr0_word_enable[31]} == 3'b001) ? wr0_data : (({wr2_word_enable[31],wr1_word_enable[31],wr0_word_enable[31]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[31],wr1_word_enable[31],wr0_word_enable[31]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1055:1024] = ({wr2_word_enable[32],wr1_word_enable[32],wr0_word_enable[32]} == 3'b001) ? wr0_data : (({wr2_word_enable[32],wr1_word_enable[32],wr0_word_enable[32]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[32],wr1_word_enable[32],wr0_word_enable[32]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1087:1056] = ({wr2_word_enable[33],wr1_word_enable[33],wr0_word_enable[33]} == 3'b001) ? wr0_data : (({wr2_word_enable[33],wr1_word_enable[33],wr0_word_enable[33]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[33],wr1_word_enable[33],wr0_word_enable[33]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1119:1088] = ({wr2_word_enable[34],wr1_word_enable[34],wr0_word_enable[34]} == 3'b001) ? wr0_data : (({wr2_word_enable[34],wr1_word_enable[34],wr0_word_enable[34]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[34],wr1_word_enable[34],wr0_word_enable[34]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1151:1120] = ({wr2_word_enable[35],wr1_word_enable[35],wr0_word_enable[35]} == 3'b001) ? wr0_data : (({wr2_word_enable[35],wr1_word_enable[35],wr0_word_enable[35]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[35],wr1_word_enable[35],wr0_word_enable[35]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1183:1152] = ({wr2_word_enable[36],wr1_word_enable[36],wr0_word_enable[36]} == 3'b001) ? wr0_data : (({wr2_word_enable[36],wr1_word_enable[36],wr0_word_enable[36]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[36],wr1_word_enable[36],wr0_word_enable[36]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1215:1184] = ({wr2_word_enable[37],wr1_word_enable[37],wr0_word_enable[37]} == 3'b001) ? wr0_data : (({wr2_word_enable[37],wr1_word_enable[37],wr0_word_enable[37]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[37],wr1_word_enable[37],wr0_word_enable[37]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1247:1216] = ({wr2_word_enable[38],wr1_word_enable[38],wr0_word_enable[38]} == 3'b001) ? wr0_data : (({wr2_word_enable[38],wr1_word_enable[38],wr0_word_enable[38]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[38],wr1_word_enable[38],wr0_word_enable[38]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1279:1248] = ({wr2_word_enable[39],wr1_word_enable[39],wr0_word_enable[39]} == 3'b001) ? wr0_data : (({wr2_word_enable[39],wr1_word_enable[39],wr0_word_enable[39]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[39],wr1_word_enable[39],wr0_word_enable[39]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1311:1280] = ({wr2_word_enable[40],wr1_word_enable[40],wr0_word_enable[40]} == 3'b001) ? wr0_data : (({wr2_word_enable[40],wr1_word_enable[40],wr0_word_enable[40]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[40],wr1_word_enable[40],wr0_word_enable[40]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1343:1312] = ({wr2_word_enable[41],wr1_word_enable[41],wr0_word_enable[41]} == 3'b001) ? wr0_data : (({wr2_word_enable[41],wr1_word_enable[41],wr0_word_enable[41]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[41],wr1_word_enable[41],wr0_word_enable[41]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1375:1344] = ({wr2_word_enable[42],wr1_word_enable[42],wr0_word_enable[42]} == 3'b001) ? wr0_data : (({wr2_word_enable[42],wr1_word_enable[42],wr0_word_enable[42]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[42],wr1_word_enable[42],wr0_word_enable[42]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1407:1376] = ({wr2_word_enable[43],wr1_word_enable[43],wr0_word_enable[43]} == 3'b001) ? wr0_data : (({wr2_word_enable[43],wr1_word_enable[43],wr0_word_enable[43]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[43],wr1_word_enable[43],wr0_word_enable[43]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1439:1408] = ({wr2_word_enable[44],wr1_word_enable[44],wr0_word_enable[44]} == 3'b001) ? wr0_data : (({wr2_word_enable[44],wr1_word_enable[44],wr0_word_enable[44]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[44],wr1_word_enable[44],wr0_word_enable[44]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1471:1440] = ({wr2_word_enable[45],wr1_word_enable[45],wr0_word_enable[45]} == 3'b001) ? wr0_data : (({wr2_word_enable[45],wr1_word_enable[45],wr0_word_enable[45]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[45],wr1_word_enable[45],wr0_word_enable[45]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1503:1472] = ({wr2_word_enable[46],wr1_word_enable[46],wr0_word_enable[46]} == 3'b001) ? wr0_data : (({wr2_word_enable[46],wr1_word_enable[46],wr0_word_enable[46]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[46],wr1_word_enable[46],wr0_word_enable[46]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1535:1504] = ({wr2_word_enable[47],wr1_word_enable[47],wr0_word_enable[47]} == 3'b001) ? wr0_data : (({wr2_word_enable[47],wr1_word_enable[47],wr0_word_enable[47]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[47],wr1_word_enable[47],wr0_word_enable[47]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1567:1536] = ({wr2_word_enable[48],wr1_word_enable[48],wr0_word_enable[48]} == 3'b001) ? wr0_data : (({wr2_word_enable[48],wr1_word_enable[48],wr0_word_enable[48]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[48],wr1_word_enable[48],wr0_word_enable[48]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1599:1568] = ({wr2_word_enable[49],wr1_word_enable[49],wr0_word_enable[49]} == 3'b001) ? wr0_data : (({wr2_word_enable[49],wr1_word_enable[49],wr0_word_enable[49]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[49],wr1_word_enable[49],wr0_word_enable[49]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1631:1600] = ({wr2_word_enable[50],wr1_word_enable[50],wr0_word_enable[50]} == 3'b001) ? wr0_data : (({wr2_word_enable[50],wr1_word_enable[50],wr0_word_enable[50]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[50],wr1_word_enable[50],wr0_word_enable[50]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1663:1632] = ({wr2_word_enable[51],wr1_word_enable[51],wr0_word_enable[51]} == 3'b001) ? wr0_data : (({wr2_word_enable[51],wr1_word_enable[51],wr0_word_enable[51]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[51],wr1_word_enable[51],wr0_word_enable[51]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1695:1664] = ({wr2_word_enable[52],wr1_word_enable[52],wr0_word_enable[52]} == 3'b001) ? wr0_data : (({wr2_word_enable[52],wr1_word_enable[52],wr0_word_enable[52]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[52],wr1_word_enable[52],wr0_word_enable[52]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1727:1696] = ({wr2_word_enable[53],wr1_word_enable[53],wr0_word_enable[53]} == 3'b001) ? wr0_data : (({wr2_word_enable[53],wr1_word_enable[53],wr0_word_enable[53]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[53],wr1_word_enable[53],wr0_word_enable[53]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1759:1728] = ({wr2_word_enable[54],wr1_word_enable[54],wr0_word_enable[54]} == 3'b001) ? wr0_data : (({wr2_word_enable[54],wr1_word_enable[54],wr0_word_enable[54]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[54],wr1_word_enable[54],wr0_word_enable[54]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1791:1760] = ({wr2_word_enable[55],wr1_word_enable[55],wr0_word_enable[55]} == 3'b001) ? wr0_data : (({wr2_word_enable[55],wr1_word_enable[55],wr0_word_enable[55]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[55],wr1_word_enable[55],wr0_word_enable[55]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1823:1792] = ({wr2_word_enable[56],wr1_word_enable[56],wr0_word_enable[56]} == 3'b001) ? wr0_data : (({wr2_word_enable[56],wr1_word_enable[56],wr0_word_enable[56]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[56],wr1_word_enable[56],wr0_word_enable[56]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1855:1824] = ({wr2_word_enable[57],wr1_word_enable[57],wr0_word_enable[57]} == 3'b001) ? wr0_data : (({wr2_word_enable[57],wr1_word_enable[57],wr0_word_enable[57]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[57],wr1_word_enable[57],wr0_word_enable[57]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1887:1856] = ({wr2_word_enable[58],wr1_word_enable[58],wr0_word_enable[58]} == 3'b001) ? wr0_data : (({wr2_word_enable[58],wr1_word_enable[58],wr0_word_enable[58]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[58],wr1_word_enable[58],wr0_word_enable[58]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1919:1888] = ({wr2_word_enable[59],wr1_word_enable[59],wr0_word_enable[59]} == 3'b001) ? wr0_data : (({wr2_word_enable[59],wr1_word_enable[59],wr0_word_enable[59]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[59],wr1_word_enable[59],wr0_word_enable[59]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1951:1920] = ({wr2_word_enable[60],wr1_word_enable[60],wr0_word_enable[60]} == 3'b001) ? wr0_data : (({wr2_word_enable[60],wr1_word_enable[60],wr0_word_enable[60]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[60],wr1_word_enable[60],wr0_word_enable[60]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[1983:1952] = ({wr2_word_enable[61],wr1_word_enable[61],wr0_word_enable[61]} == 3'b001) ? wr0_data : (({wr2_word_enable[61],wr1_word_enable[61],wr0_word_enable[61]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[61],wr1_word_enable[61],wr0_word_enable[61]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2015:1984] = ({wr2_word_enable[62],wr1_word_enable[62],wr0_word_enable[62]} == 3'b001) ? wr0_data : (({wr2_word_enable[62],wr1_word_enable[62],wr0_word_enable[62]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[62],wr1_word_enable[62],wr0_word_enable[62]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2047:2016] = ({wr2_word_enable[63],wr1_word_enable[63],wr0_word_enable[63]} == 3'b001) ? wr0_data : (({wr2_word_enable[63],wr1_word_enable[63],wr0_word_enable[63]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[63],wr1_word_enable[63],wr0_word_enable[63]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2079:2048] = ({wr2_word_enable[64],wr1_word_enable[64],wr0_word_enable[64]} == 3'b001) ? wr0_data : (({wr2_word_enable[64],wr1_word_enable[64],wr0_word_enable[64]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[64],wr1_word_enable[64],wr0_word_enable[64]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2111:2080] = ({wr2_word_enable[65],wr1_word_enable[65],wr0_word_enable[65]} == 3'b001) ? wr0_data : (({wr2_word_enable[65],wr1_word_enable[65],wr0_word_enable[65]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[65],wr1_word_enable[65],wr0_word_enable[65]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2143:2112] = ({wr2_word_enable[66],wr1_word_enable[66],wr0_word_enable[66]} == 3'b001) ? wr0_data : (({wr2_word_enable[66],wr1_word_enable[66],wr0_word_enable[66]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[66],wr1_word_enable[66],wr0_word_enable[66]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2175:2144] = ({wr2_word_enable[67],wr1_word_enable[67],wr0_word_enable[67]} == 3'b001) ? wr0_data : (({wr2_word_enable[67],wr1_word_enable[67],wr0_word_enable[67]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[67],wr1_word_enable[67],wr0_word_enable[67]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2207:2176] = ({wr2_word_enable[68],wr1_word_enable[68],wr0_word_enable[68]} == 3'b001) ? wr0_data : (({wr2_word_enable[68],wr1_word_enable[68],wr0_word_enable[68]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[68],wr1_word_enable[68],wr0_word_enable[68]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2239:2208] = ({wr2_word_enable[69],wr1_word_enable[69],wr0_word_enable[69]} == 3'b001) ? wr0_data : (({wr2_word_enable[69],wr1_word_enable[69],wr0_word_enable[69]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[69],wr1_word_enable[69],wr0_word_enable[69]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2271:2240] = ({wr2_word_enable[70],wr1_word_enable[70],wr0_word_enable[70]} == 3'b001) ? wr0_data : (({wr2_word_enable[70],wr1_word_enable[70],wr0_word_enable[70]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[70],wr1_word_enable[70],wr0_word_enable[70]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2303:2272] = ({wr2_word_enable[71],wr1_word_enable[71],wr0_word_enable[71]} == 3'b001) ? wr0_data : (({wr2_word_enable[71],wr1_word_enable[71],wr0_word_enable[71]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[71],wr1_word_enable[71],wr0_word_enable[71]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2335:2304] = ({wr2_word_enable[72],wr1_word_enable[72],wr0_word_enable[72]} == 3'b001) ? wr0_data : (({wr2_word_enable[72],wr1_word_enable[72],wr0_word_enable[72]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[72],wr1_word_enable[72],wr0_word_enable[72]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2367:2336] = ({wr2_word_enable[73],wr1_word_enable[73],wr0_word_enable[73]} == 3'b001) ? wr0_data : (({wr2_word_enable[73],wr1_word_enable[73],wr0_word_enable[73]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[73],wr1_word_enable[73],wr0_word_enable[73]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2399:2368] = ({wr2_word_enable[74],wr1_word_enable[74],wr0_word_enable[74]} == 3'b001) ? wr0_data : (({wr2_word_enable[74],wr1_word_enable[74],wr0_word_enable[74]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[74],wr1_word_enable[74],wr0_word_enable[74]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2431:2400] = ({wr2_word_enable[75],wr1_word_enable[75],wr0_word_enable[75]} == 3'b001) ? wr0_data : (({wr2_word_enable[75],wr1_word_enable[75],wr0_word_enable[75]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[75],wr1_word_enable[75],wr0_word_enable[75]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2463:2432] = ({wr2_word_enable[76],wr1_word_enable[76],wr0_word_enable[76]} == 3'b001) ? wr0_data : (({wr2_word_enable[76],wr1_word_enable[76],wr0_word_enable[76]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[76],wr1_word_enable[76],wr0_word_enable[76]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2495:2464] = ({wr2_word_enable[77],wr1_word_enable[77],wr0_word_enable[77]} == 3'b001) ? wr0_data : (({wr2_word_enable[77],wr1_word_enable[77],wr0_word_enable[77]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[77],wr1_word_enable[77],wr0_word_enable[77]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2527:2496] = ({wr2_word_enable[78],wr1_word_enable[78],wr0_word_enable[78]} == 3'b001) ? wr0_data : (({wr2_word_enable[78],wr1_word_enable[78],wr0_word_enable[78]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[78],wr1_word_enable[78],wr0_word_enable[78]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2559:2528] = ({wr2_word_enable[79],wr1_word_enable[79],wr0_word_enable[79]} == 3'b001) ? wr0_data : (({wr2_word_enable[79],wr1_word_enable[79],wr0_word_enable[79]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[79],wr1_word_enable[79],wr0_word_enable[79]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2591:2560] = ({wr2_word_enable[80],wr1_word_enable[80],wr0_word_enable[80]} == 3'b001) ? wr0_data : (({wr2_word_enable[80],wr1_word_enable[80],wr0_word_enable[80]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[80],wr1_word_enable[80],wr0_word_enable[80]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2623:2592] = ({wr2_word_enable[81],wr1_word_enable[81],wr0_word_enable[81]} == 3'b001) ? wr0_data : (({wr2_word_enable[81],wr1_word_enable[81],wr0_word_enable[81]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[81],wr1_word_enable[81],wr0_word_enable[81]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2655:2624] = ({wr2_word_enable[82],wr1_word_enable[82],wr0_word_enable[82]} == 3'b001) ? wr0_data : (({wr2_word_enable[82],wr1_word_enable[82],wr0_word_enable[82]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[82],wr1_word_enable[82],wr0_word_enable[82]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2687:2656] = ({wr2_word_enable[83],wr1_word_enable[83],wr0_word_enable[83]} == 3'b001) ? wr0_data : (({wr2_word_enable[83],wr1_word_enable[83],wr0_word_enable[83]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[83],wr1_word_enable[83],wr0_word_enable[83]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2719:2688] = ({wr2_word_enable[84],wr1_word_enable[84],wr0_word_enable[84]} == 3'b001) ? wr0_data : (({wr2_word_enable[84],wr1_word_enable[84],wr0_word_enable[84]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[84],wr1_word_enable[84],wr0_word_enable[84]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2751:2720] = ({wr2_word_enable[85],wr1_word_enable[85],wr0_word_enable[85]} == 3'b001) ? wr0_data : (({wr2_word_enable[85],wr1_word_enable[85],wr0_word_enable[85]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[85],wr1_word_enable[85],wr0_word_enable[85]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2783:2752] = ({wr2_word_enable[86],wr1_word_enable[86],wr0_word_enable[86]} == 3'b001) ? wr0_data : (({wr2_word_enable[86],wr1_word_enable[86],wr0_word_enable[86]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[86],wr1_word_enable[86],wr0_word_enable[86]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2815:2784] = ({wr2_word_enable[87],wr1_word_enable[87],wr0_word_enable[87]} == 3'b001) ? wr0_data : (({wr2_word_enable[87],wr1_word_enable[87],wr0_word_enable[87]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[87],wr1_word_enable[87],wr0_word_enable[87]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2847:2816] = ({wr2_word_enable[88],wr1_word_enable[88],wr0_word_enable[88]} == 3'b001) ? wr0_data : (({wr2_word_enable[88],wr1_word_enable[88],wr0_word_enable[88]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[88],wr1_word_enable[88],wr0_word_enable[88]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2879:2848] = ({wr2_word_enable[89],wr1_word_enable[89],wr0_word_enable[89]} == 3'b001) ? wr0_data : (({wr2_word_enable[89],wr1_word_enable[89],wr0_word_enable[89]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[89],wr1_word_enable[89],wr0_word_enable[89]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2911:2880] = ({wr2_word_enable[90],wr1_word_enable[90],wr0_word_enable[90]} == 3'b001) ? wr0_data : (({wr2_word_enable[90],wr1_word_enable[90],wr0_word_enable[90]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[90],wr1_word_enable[90],wr0_word_enable[90]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2943:2912] = ({wr2_word_enable[91],wr1_word_enable[91],wr0_word_enable[91]} == 3'b001) ? wr0_data : (({wr2_word_enable[91],wr1_word_enable[91],wr0_word_enable[91]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[91],wr1_word_enable[91],wr0_word_enable[91]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[2975:2944] = ({wr2_word_enable[92],wr1_word_enable[92],wr0_word_enable[92]} == 3'b001) ? wr0_data : (({wr2_word_enable[92],wr1_word_enable[92],wr0_word_enable[92]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[92],wr1_word_enable[92],wr0_word_enable[92]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3007:2976] = ({wr2_word_enable[93],wr1_word_enable[93],wr0_word_enable[93]} == 3'b001) ? wr0_data : (({wr2_word_enable[93],wr1_word_enable[93],wr0_word_enable[93]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[93],wr1_word_enable[93],wr0_word_enable[93]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3039:3008] = ({wr2_word_enable[94],wr1_word_enable[94],wr0_word_enable[94]} == 3'b001) ? wr0_data : (({wr2_word_enable[94],wr1_word_enable[94],wr0_word_enable[94]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[94],wr1_word_enable[94],wr0_word_enable[94]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3071:3040] = ({wr2_word_enable[95],wr1_word_enable[95],wr0_word_enable[95]} == 3'b001) ? wr0_data : (({wr2_word_enable[95],wr1_word_enable[95],wr0_word_enable[95]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[95],wr1_word_enable[95],wr0_word_enable[95]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3103:3072] = ({wr2_word_enable[96],wr1_word_enable[96],wr0_word_enable[96]} == 3'b001) ? wr0_data : (({wr2_word_enable[96],wr1_word_enable[96],wr0_word_enable[96]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[96],wr1_word_enable[96],wr0_word_enable[96]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3135:3104] = ({wr2_word_enable[97],wr1_word_enable[97],wr0_word_enable[97]} == 3'b001) ? wr0_data : (({wr2_word_enable[97],wr1_word_enable[97],wr0_word_enable[97]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[97],wr1_word_enable[97],wr0_word_enable[97]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3167:3136] = ({wr2_word_enable[98],wr1_word_enable[98],wr0_word_enable[98]} == 3'b001) ? wr0_data : (({wr2_word_enable[98],wr1_word_enable[98],wr0_word_enable[98]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[98],wr1_word_enable[98],wr0_word_enable[98]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3199:3168] = ({wr2_word_enable[99],wr1_word_enable[99],wr0_word_enable[99]} == 3'b001) ? wr0_data : (({wr2_word_enable[99],wr1_word_enable[99],wr0_word_enable[99]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[99],wr1_word_enable[99],wr0_word_enable[99]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3231:3200] = ({wr2_word_enable[100],wr1_word_enable[100],wr0_word_enable[100]} == 3'b001) ? wr0_data : (({wr2_word_enable[100],wr1_word_enable[100],wr0_word_enable[100]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[100],wr1_word_enable[100],wr0_word_enable[100]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3263:3232] = ({wr2_word_enable[101],wr1_word_enable[101],wr0_word_enable[101]} == 3'b001) ? wr0_data : (({wr2_word_enable[101],wr1_word_enable[101],wr0_word_enable[101]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[101],wr1_word_enable[101],wr0_word_enable[101]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3295:3264] = ({wr2_word_enable[102],wr1_word_enable[102],wr0_word_enable[102]} == 3'b001) ? wr0_data : (({wr2_word_enable[102],wr1_word_enable[102],wr0_word_enable[102]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[102],wr1_word_enable[102],wr0_word_enable[102]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3327:3296] = ({wr2_word_enable[103],wr1_word_enable[103],wr0_word_enable[103]} == 3'b001) ? wr0_data : (({wr2_word_enable[103],wr1_word_enable[103],wr0_word_enable[103]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[103],wr1_word_enable[103],wr0_word_enable[103]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3359:3328] = ({wr2_word_enable[104],wr1_word_enable[104],wr0_word_enable[104]} == 3'b001) ? wr0_data : (({wr2_word_enable[104],wr1_word_enable[104],wr0_word_enable[104]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[104],wr1_word_enable[104],wr0_word_enable[104]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3391:3360] = ({wr2_word_enable[105],wr1_word_enable[105],wr0_word_enable[105]} == 3'b001) ? wr0_data : (({wr2_word_enable[105],wr1_word_enable[105],wr0_word_enable[105]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[105],wr1_word_enable[105],wr0_word_enable[105]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3423:3392] = ({wr2_word_enable[106],wr1_word_enable[106],wr0_word_enable[106]} == 3'b001) ? wr0_data : (({wr2_word_enable[106],wr1_word_enable[106],wr0_word_enable[106]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[106],wr1_word_enable[106],wr0_word_enable[106]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3455:3424] = ({wr2_word_enable[107],wr1_word_enable[107],wr0_word_enable[107]} == 3'b001) ? wr0_data : (({wr2_word_enable[107],wr1_word_enable[107],wr0_word_enable[107]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[107],wr1_word_enable[107],wr0_word_enable[107]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3487:3456] = ({wr2_word_enable[108],wr1_word_enable[108],wr0_word_enable[108]} == 3'b001) ? wr0_data : (({wr2_word_enable[108],wr1_word_enable[108],wr0_word_enable[108]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[108],wr1_word_enable[108],wr0_word_enable[108]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3519:3488] = ({wr2_word_enable[109],wr1_word_enable[109],wr0_word_enable[109]} == 3'b001) ? wr0_data : (({wr2_word_enable[109],wr1_word_enable[109],wr0_word_enable[109]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[109],wr1_word_enable[109],wr0_word_enable[109]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3551:3520] = ({wr2_word_enable[110],wr1_word_enable[110],wr0_word_enable[110]} == 3'b001) ? wr0_data : (({wr2_word_enable[110],wr1_word_enable[110],wr0_word_enable[110]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[110],wr1_word_enable[110],wr0_word_enable[110]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3583:3552] = ({wr2_word_enable[111],wr1_word_enable[111],wr0_word_enable[111]} == 3'b001) ? wr0_data : (({wr2_word_enable[111],wr1_word_enable[111],wr0_word_enable[111]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[111],wr1_word_enable[111],wr0_word_enable[111]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3615:3584] = ({wr2_word_enable[112],wr1_word_enable[112],wr0_word_enable[112]} == 3'b001) ? wr0_data : (({wr2_word_enable[112],wr1_word_enable[112],wr0_word_enable[112]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[112],wr1_word_enable[112],wr0_word_enable[112]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3647:3616] = ({wr2_word_enable[113],wr1_word_enable[113],wr0_word_enable[113]} == 3'b001) ? wr0_data : (({wr2_word_enable[113],wr1_word_enable[113],wr0_word_enable[113]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[113],wr1_word_enable[113],wr0_word_enable[113]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3679:3648] = ({wr2_word_enable[114],wr1_word_enable[114],wr0_word_enable[114]} == 3'b001) ? wr0_data : (({wr2_word_enable[114],wr1_word_enable[114],wr0_word_enable[114]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[114],wr1_word_enable[114],wr0_word_enable[114]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3711:3680] = ({wr2_word_enable[115],wr1_word_enable[115],wr0_word_enable[115]} == 3'b001) ? wr0_data : (({wr2_word_enable[115],wr1_word_enable[115],wr0_word_enable[115]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[115],wr1_word_enable[115],wr0_word_enable[115]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3743:3712] = ({wr2_word_enable[116],wr1_word_enable[116],wr0_word_enable[116]} == 3'b001) ? wr0_data : (({wr2_word_enable[116],wr1_word_enable[116],wr0_word_enable[116]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[116],wr1_word_enable[116],wr0_word_enable[116]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3775:3744] = ({wr2_word_enable[117],wr1_word_enable[117],wr0_word_enable[117]} == 3'b001) ? wr0_data : (({wr2_word_enable[117],wr1_word_enable[117],wr0_word_enable[117]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[117],wr1_word_enable[117],wr0_word_enable[117]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3807:3776] = ({wr2_word_enable[118],wr1_word_enable[118],wr0_word_enable[118]} == 3'b001) ? wr0_data : (({wr2_word_enable[118],wr1_word_enable[118],wr0_word_enable[118]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[118],wr1_word_enable[118],wr0_word_enable[118]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3839:3808] = ({wr2_word_enable[119],wr1_word_enable[119],wr0_word_enable[119]} == 3'b001) ? wr0_data : (({wr2_word_enable[119],wr1_word_enable[119],wr0_word_enable[119]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[119],wr1_word_enable[119],wr0_word_enable[119]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3871:3840] = ({wr2_word_enable[120],wr1_word_enable[120],wr0_word_enable[120]} == 3'b001) ? wr0_data : (({wr2_word_enable[120],wr1_word_enable[120],wr0_word_enable[120]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[120],wr1_word_enable[120],wr0_word_enable[120]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3903:3872] = ({wr2_word_enable[121],wr1_word_enable[121],wr0_word_enable[121]} == 3'b001) ? wr0_data : (({wr2_word_enable[121],wr1_word_enable[121],wr0_word_enable[121]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[121],wr1_word_enable[121],wr0_word_enable[121]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3935:3904] = ({wr2_word_enable[122],wr1_word_enable[122],wr0_word_enable[122]} == 3'b001) ? wr0_data : (({wr2_word_enable[122],wr1_word_enable[122],wr0_word_enable[122]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[122],wr1_word_enable[122],wr0_word_enable[122]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3967:3936] = ({wr2_word_enable[123],wr1_word_enable[123],wr0_word_enable[123]} == 3'b001) ? wr0_data : (({wr2_word_enable[123],wr1_word_enable[123],wr0_word_enable[123]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[123],wr1_word_enable[123],wr0_word_enable[123]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[3999:3968] = ({wr2_word_enable[124],wr1_word_enable[124],wr0_word_enable[124]} == 3'b001) ? wr0_data : (({wr2_word_enable[124],wr1_word_enable[124],wr0_word_enable[124]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[124],wr1_word_enable[124],wr0_word_enable[124]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[4031:4000] = ({wr2_word_enable[125],wr1_word_enable[125],wr0_word_enable[125]} == 3'b001) ? wr0_data : (({wr2_word_enable[125],wr1_word_enable[125],wr0_word_enable[125]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[125],wr1_word_enable[125],wr0_word_enable[125]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[4063:4032] = ({wr2_word_enable[126],wr1_word_enable[126],wr0_word_enable[126]} == 3'b001) ? wr0_data : (({wr2_word_enable[126],wr1_word_enable[126],wr0_word_enable[126]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[126],wr1_word_enable[126],wr0_word_enable[126]} == 3'b100)? wr2_data : {32{1'bx}}));
assign word_in[4095:4064] = ({wr2_word_enable[127],wr1_word_enable[127],wr0_word_enable[127]} == 3'b001) ? wr0_data : (({wr2_word_enable[127],wr1_word_enable[127],wr0_word_enable[127]} == 3'b010) ? wr1_data : ( ({wr2_word_enable[127],wr1_word_enable[127],wr0_word_enable[127]} == 3'b100)? wr2_data : {32{1'bx}}));

endmodule
